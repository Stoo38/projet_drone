../../BENCH/tbench.sv