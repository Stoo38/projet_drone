../results/top_ppm.vhd