../../BENCH/tbench_sans_top.sv