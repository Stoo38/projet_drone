../results/top_bar.vhd