../../BENCH/test_counter.vhd