
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_bar is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_top_bar;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_bar.all;

entity top_bar is

   port( CLK_top, reset_top, SW1_top : in std_logic;  r_top, g_top, b_top : in 
         std_logic_vector (7 downto 0);  rout_top, gout_top, bout_top, 
         r_out_proc, g_out_proc, b_out_proc : out std_logic_vector (7 downto 0)
         ;  X_barycentre_top, Y_barycentre_top : out std_logic_vector (8 downto
         0);  HSYNC_top, VSYNC_top : out std_logic;  cam_x : out 
         std_logic_vector (9 downto 0);  cam_y : out std_logic_vector (8 downto
         0);  IMG_top : out std_logic);

end top_bar;

architecture SYN_bar of top_bar is

   component OAI212
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI222
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component IMAJ31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component LOGIC1
      port( Q : out std_logic);
   end component;
   
   component BUF2
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component INV3
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR40
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI221
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND22
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI211
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR41
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI311
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND41
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI311
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component BUF6
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component MAJ31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component DFE1
      port( D, E, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component DF3
      port( D, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLPQ3
      port( SN, D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component ADD22
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADD32
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal r_out_proc_7_port, r_out_proc_6_port, r_out_proc_5_port, 
      r_out_proc_4_port, r_out_proc_3_port, r_out_proc_2_port, 
      r_out_proc_1_port, r_out_proc_0_port, g_out_proc_7_port, 
      g_out_proc_6_port, g_out_proc_5_port, g_out_proc_4_port, 
      g_out_proc_3_port, g_out_proc_2_port, g_out_proc_1_port, 
      g_out_proc_0_port, b_out_proc_7_port, b_out_proc_6_port, 
      b_out_proc_5_port, b_out_proc_4_port, b_out_proc_3_port, 
      b_out_proc_2_port, b_out_proc_1_port, b_out_proc_0_port, 
      X_barycentre_top_8_port, X_barycentre_top_7_port, X_barycentre_top_6_port
      , X_barycentre_top_5_port, X_barycentre_top_4_port, 
      X_barycentre_top_3_port, X_barycentre_top_2_port, X_barycentre_top_1_port
      , X_barycentre_top_0_port, Y_barycentre_top_8_port, 
      Y_barycentre_top_7_port, Y_barycentre_top_6_port, Y_barycentre_top_5_port
      , Y_barycentre_top_4_port, Y_barycentre_top_3_port, 
      Y_barycentre_top_2_port, Y_barycentre_top_1_port, Y_barycentre_top_0_port
      , cam_x_9_port, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, 
      n2136, gensync1_n107, gensync1_n106, gensync1_n105, gensync1_n104, 
      gensync1_n103, gensync1_n102, gensync1_n101, gensync1_n100, gensync1_n99,
      gensync1_n98, gensync1_n97, gensync1_n96, gensync1_n95, gensync1_n94, 
      gensync1_n93, gensync1_n92, gensync1_n91, gensync1_n90, gensync1_n89, 
      gensync1_n88, gensync1_n87, gensync1_N182, gensync1_N181, gensync1_N180, 
      gensync1_N179, gensync1_N178, gensync1_N177, gensync1_N176, gensync1_N175
      , gensync1_N174, gensync1_N173, gensync1_N172, gensync1_N171, 
      gensync1_N170, gensync1_N169, gensync1_N168, gensync1_N167, gensync1_N166
      , gensync1_N165, gensync1_N145, gensync1_N144, gensync1_N143, 
      gensync1_N142, gensync1_N141, gensync1_N140, gensync1_N139, gensync1_N138
      , gensync1_N135, gensync1_N132, gensync1_N129, gensync1_N85, gensync1_N74
      , gensync1_N72, gensync1_N69, gensync1_N66, gensync1_N65, gensync1_N64, 
      gensync1_N63, gensync1_N62, gensync1_N61, gensync1_N60, gensync1_N59, 
      gensync1_N58, gensync1_N57, gensync1_N56, gensync1_N54, gensync1_N53, 
      gensync1_N52, gensync1_N51, gensync1_N50, gensync1_N49, gensync1_N48, 
      gensync1_N47, gensync1_N43, gensync1_comptY_9_port, gensync1_N31, 
      gensync1_N30, gensync1_N29, gensync1_N28, gensync1_N27, gensync1_N26, 
      gensync1_N25, gensync1_N24, gensync1_N23, gensync1_N22, gensync1_N20, 
      gensync1_N19, gensync1_N18, gensync1_N17, gensync1_N16, gensync1_N15, 
      gensync1_N14, gensync1_N13, gensync1_N9, image_process1_n119, 
      image_process1_n118, image_process1_n117, image_process1_n116, 
      image_process1_n115, image_process1_n114, image_process1_n113, 
      image_process1_n112, image_process1_n111, image_process1_n110, 
      image_process1_n109, image_process1_n108, image_process1_n107, 
      image_process1_n106, image_process1_n105, image_process1_n104, 
      image_process1_n103, image_process1_n102, image_process1_n101, 
      image_process1_n100, image_process1_n99, image_process1_n98, 
      image_process1_n97, image_process1_n96, image_process1_n95, 
      image_process1_n94, image_process1_n93, image_process1_n92, 
      image_process1_n91, image_process1_n90, image_process1_n89, 
      image_process1_n88, image_process1_n87, image_process1_n86, 
      image_process1_n85, image_process1_n84, image_process1_n83, 
      image_process1_n82, image_process1_n81, image_process1_n80, 
      image_process1_n79, image_process1_n78, image_process1_n77, 
      image_process1_n76, image_process1_n75, image_process1_n74, 
      image_process1_n73, image_process1_n72, image_process1_n71, 
      image_process1_n70, image_process1_n69, image_process1_n68, 
      image_process1_n67, image_process1_n66, image_process1_n65, 
      image_process1_n64, image_process1_n63, image_process1_n62, 
      image_process1_n61, image_process1_n60, image_process1_n59, 
      image_process1_n58, image_process1_n57, image_process1_n56, 
      image_process1_n55, image_process1_n27, image_process1_n25, 
      image_process1_n13, image_process1_N64_port, image_process1_N62_port, 
      image_process1_N59_port, image_process1_N31, image_process1_N29, 
      image_process1_N28, image_process1_N26, image_process1_N25_port, 
      image_process1_N23, image_process1_N22, image_process1_N20, 
      image_process1_N19, image_process1_N17, image_process1_N16, 
      image_process1_N14, image_process1_N13_port, image_process1_N11, 
      image_process1_N10, image_process1_N8, image_process1_state, 
      image_process1_bi_0_port, image_process1_bi_1_port, 
      image_process1_bi_3_port, image_process1_bi_4_port, 
      image_process1_bi_5_port, image_process1_bi_6_port, 
      image_process1_bi_7_port, image_process1_gi_0_port, 
      image_process1_gi_1_port, image_process1_gi_2_port, 
      image_process1_gi_3_port, image_process1_gi_4_port, 
      image_process1_gi_5_port, image_process1_gi_6_port, 
      image_process1_gi_7_port, image_process1_ri_0_port, 
      image_process1_ri_1_port, image_process1_ri_3_port, 
      image_process1_ri_4_port, image_process1_ri_5_port, 
      image_process1_ri_6_port, image_process1_ri_7_port, position1_n1635, 
      position1_n1634, position1_n1633, position1_n1632, position1_n1631, 
      position1_n1630, position1_n1629, position1_n1628, position1_n1627, 
      position1_n1626, position1_n1625, position1_n1624, position1_n1623, 
      position1_n1622, position1_n1621, position1_n1620, position1_n1619, 
      position1_n1618, position1_n1617, position1_n1616, position1_n1615, 
      position1_n1614, position1_n1613, position1_n1612, position1_n1611, 
      position1_n1610, position1_n1609, position1_n1608, position1_n1607, 
      position1_n1606, position1_n1605, position1_n1604, position1_n1603, 
      position1_n1602, position1_n1601, position1_n1600, position1_n1599, 
      position1_n1598, position1_n1597, position1_n1596, position1_n1595, 
      position1_n1594, position1_n1593, position1_n1592, position1_n1591, 
      position1_n1590, position1_n1589, position1_n1588, position1_n1587, 
      position1_n1586, position1_n1585, position1_n1584, position1_n1583, 
      position1_n1582, position1_n1581, position1_n1580, position1_n1579, 
      position1_n1578, position1_n1577, position1_n1576, position1_n1575, 
      position1_n1574, position1_n1573, position1_n1572, position1_n1571, 
      position1_n1570, position1_n1569, position1_n1568, position1_n1567, 
      position1_n1566, position1_n1565, position1_n1564, position1_n1563, 
      position1_n1562, position1_n1561, position1_n1560, position1_n1559, 
      position1_n1558, position1_n1557, position1_n1556, position1_n1555, 
      position1_n1554, position1_n1553, position1_n1552, position1_n1551, 
      position1_n1550, position1_n1549, position1_n1548, position1_n1547, 
      position1_n1546, position1_n1545, position1_n1544, position1_n1543, 
      position1_n1542, position1_n1541, position1_n1540, position1_n1539, 
      position1_n1538, position1_n1537, position1_n1536, position1_n1535, 
      position1_n1534, position1_n1533, position1_n1532, position1_n1531, 
      position1_n1530, position1_n1529, position1_n1528, position1_n1527, 
      position1_n1526, position1_n1525, position1_n1524, position1_n1523, 
      position1_n1522, position1_n1521, position1_n1520, position1_n1519, 
      position1_n1518, position1_n1517, position1_n1516, position1_n1515, 
      position1_n1514, position1_n1513, position1_n1512, position1_n1511, 
      position1_n1510, position1_n1509, position1_n1508, position1_n1507, 
      position1_n1506, position1_n1505, position1_n1504, position1_n1503, 
      position1_n1502, position1_n1501, position1_n1500, position1_n1499, 
      position1_n1498, position1_n1497, position1_n1496, position1_n1495, 
      position1_n1494, position1_n1493, position1_n1492, position1_n1491, 
      position1_n1490, position1_n1489, position1_n1488, position1_n1487, 
      position1_n1486, position1_n1485, position1_n1484, position1_n1483, 
      position1_n1482, position1_n1481, position1_n1480, position1_n1479, 
      position1_n1478, position1_n1477, position1_n1476, position1_n1475, 
      position1_n1474, position1_n1473, position1_n1472, position1_n1471, 
      position1_n1470, position1_n1469, position1_n1468, position1_n1467, 
      position1_n1466, position1_n1465, position1_n1464, position1_n1463, 
      position1_n1462, position1_n1461, position1_n1460, position1_n1459, 
      position1_n1458, position1_n1457, position1_n1456, position1_n1455, 
      position1_n1454, position1_n1453, position1_n1452, position1_n1451, 
      position1_n1450, position1_n1449, position1_n1448, position1_n1447, 
      position1_n1446, position1_n1445, position1_n1444, position1_n1443, 
      position1_n1442, position1_n1441, position1_n1440, position1_n1439, 
      position1_n1438, position1_n1437, position1_n1436, position1_n1435, 
      position1_n1434, position1_n1433, position1_n1432, position1_n1431, 
      position1_n1430, position1_n1429, position1_n1428, position1_n1427, 
      position1_n1426, position1_n1425, position1_n1424, position1_n1423, 
      position1_n1422, position1_n1421, position1_n1420, position1_n1419, 
      position1_n1418, position1_n1417, position1_n1416, position1_n1415, 
      position1_n1414, position1_n1413, position1_n1412, position1_n1411, 
      position1_n1410, position1_n1409, position1_n1408, position1_n1407, 
      position1_n1406, position1_n1405, position1_n1404, position1_n1403, 
      position1_n1402, position1_n1401, position1_n1400, position1_n1399, 
      position1_n1398, position1_n1397, position1_n1396, position1_n1395, 
      position1_n1394, position1_n1393, position1_n1392, position1_n1391, 
      position1_n1390, position1_n1389, position1_n1388, position1_n1387, 
      position1_n1386, position1_n1385, position1_n1384, position1_n1383, 
      position1_n1382, position1_n1381, position1_n1380, position1_n1379, 
      position1_n1378, position1_n1377, position1_n1376, position1_n1375, 
      position1_n1374, position1_n1373, position1_n1372, position1_n1371, 
      position1_n1370, position1_n1369, position1_n1368, position1_n1367, 
      position1_n1366, position1_n1365, position1_n1364, position1_n1363, 
      position1_n1362, position1_n1361, position1_n1360, position1_n1359, 
      position1_n1358, position1_n1357, position1_n1356, position1_n1355, 
      position1_n1354, position1_n1353, position1_n1352, position1_n1351, 
      position1_n1350, position1_n1349, position1_n1348, position1_n1347, 
      position1_n1346, position1_n1345, position1_n1344, position1_n1343, 
      position1_n1342, position1_n1341, position1_n1340, position1_n1339, 
      position1_n1338, position1_n1337, position1_n1336, position1_n1335, 
      position1_n1334, position1_n1333, position1_n1332, position1_n1331, 
      position1_n1330, position1_n1329, position1_n1328, position1_n1327, 
      position1_n1326, position1_n1325, position1_n1324, position1_n1323, 
      position1_n1322, position1_n1321, position1_n1320, position1_n1319, 
      position1_n1318, position1_n1317, position1_n1316, position1_n1315, 
      position1_n1314, position1_n1313, position1_n1312, position1_n1311, 
      position1_n1310, position1_n1309, position1_n1308, position1_n1307, 
      position1_n1306, position1_n1305, position1_n1304, position1_n1303, 
      position1_n1302, position1_n1301, position1_n1300, position1_n1299, 
      position1_n1298, position1_n1297, position1_n1296, position1_n1295, 
      position1_n1294, position1_n1293, position1_n1292, position1_n1291, 
      position1_n1290, position1_n1289, position1_n1288, position1_n1287, 
      position1_n1286, position1_n1285, position1_n1284, position1_n1283, 
      position1_n1282, position1_n1281, position1_n1280, position1_n1279, 
      position1_n1278, position1_n1277, position1_n1276, position1_n1275, 
      position1_n1274, position1_n1273, position1_n1272, position1_n1271, 
      position1_n1270, position1_n1269, position1_n1268, position1_n1267, 
      position1_n1266, position1_n1265, position1_n1264, position1_n1263, 
      position1_n1262, position1_n1261, position1_n1260, position1_n1259, 
      position1_n1258, position1_n1257, position1_n1256, position1_n1255, 
      position1_n1254, position1_n1253, position1_n1252, position1_n1251, 
      position1_n1250, position1_n1249, position1_n1248, position1_n1247, 
      position1_n1246, position1_n1245, position1_n1244, position1_n1243, 
      position1_n1242, position1_n1241, position1_n1240, position1_n1239, 
      position1_n1238, position1_n1237, position1_n1236, position1_n1235, 
      position1_n1234, position1_n1233, position1_n1232, position1_n1231, 
      position1_n1230, position1_n1229, position1_n1228, position1_n1227, 
      position1_n1226, position1_n1225, position1_n1224, position1_n1223, 
      position1_n1222, position1_n1221, position1_n1220, position1_n1219, 
      position1_n1218, position1_n1217, position1_n1216, position1_n1215, 
      position1_n1214, position1_n1213, position1_n1212, position1_n1211, 
      position1_n1210, position1_n1209, position1_n1208, position1_n1207, 
      position1_n1206, position1_n1205, position1_n1204, position1_n1203, 
      position1_n1202, position1_n1201, position1_n1200, position1_n1199, 
      position1_n1198, position1_n1197, position1_n1196, position1_n1195, 
      position1_n1194, position1_n1193, position1_n1192, position1_n1191, 
      position1_n1190, position1_n1189, position1_n1188, position1_n1187, 
      position1_n1186, position1_n1185, position1_n1184, position1_n1183, 
      position1_n1182, position1_n1181, position1_n1180, position1_n1179, 
      position1_n1178, position1_n1177, position1_n1176, position1_n1175, 
      position1_n1174, position1_n1173, position1_n1172, position1_n1171, 
      position1_n1170, position1_n1169, position1_n1168, position1_n1167, 
      position1_n1166, position1_n1165, position1_n1164, position1_n1163, 
      position1_n1162, position1_n1161, position1_n1160, position1_n1159, 
      position1_n1158, position1_n1157, position1_n1156, position1_n1154, 
      position1_n1153, position1_n1152, position1_n1151, position1_n1150, 
      position1_n1149, position1_n1148, position1_n1147, position1_n1146, 
      position1_n1145, position1_n1144, position1_n1143, position1_n1142, 
      position1_n1141, position1_n1140, position1_n1139, position1_n1138, 
      position1_n1137, position1_n1136, position1_n1135, position1_n1134, 
      position1_n1133, position1_n1132, position1_n1131, position1_n1130, 
      position1_n1129, position1_n1128, position1_n1127, position1_n1126, 
      position1_n1125, position1_n1124, position1_n1123, position1_n1122, 
      position1_n1121, position1_n1120, position1_n1119, position1_n1118, 
      position1_n1117, position1_n1116, position1_n1115, position1_n1114, 
      position1_n1113, position1_n1112, position1_n1111, position1_n1110, 
      position1_n1109, position1_n1108, position1_n1107, position1_n1106, 
      position1_n1105, position1_n1104, position1_n1103, position1_n1102, 
      position1_n1101, position1_n1100, position1_n1099, position1_n1098, 
      position1_n1097, position1_n1096, position1_n1095, position1_n1094, 
      position1_n1093, position1_n1092, position1_n1091, position1_n1090, 
      position1_n1089, position1_n1088, position1_n1087, position1_n1086, 
      position1_n1085, position1_n1084, position1_n1083, position1_n1082, 
      position1_n1081, position1_n1080, position1_n1079, position1_n1078, 
      position1_n1077, position1_n1076, position1_n1075, position1_n1074, 
      position1_n1073, position1_n1072, position1_n1071, position1_n1070, 
      position1_n1069, position1_n1068, position1_n1067, position1_n1066, 
      position1_n1065, position1_n1064, position1_n1063, position1_n1062, 
      position1_n1061, position1_n1060, position1_n1059, position1_n1058, 
      position1_n1057, position1_n1056, position1_n1055, position1_n1054, 
      position1_n1053, position1_n1052, position1_n1051, position1_n1050, 
      position1_n1049, position1_n1048, position1_n1047, position1_n1046, 
      position1_n1045, position1_n1044, position1_n1043, position1_n1042, 
      position1_n1041, position1_n1040, position1_n1039, position1_n1038, 
      position1_n1037, position1_n1036, position1_n1035, position1_n1034, 
      position1_n1033, position1_n1032, position1_n1031, position1_n1030, 
      position1_n1029, position1_n1028, position1_n1027, position1_n1026, 
      position1_n1025, position1_n1024, position1_n1023, position1_n1022, 
      position1_n1021, position1_n1020, position1_n1019, position1_n1018, 
      position1_n1017, position1_n1016, position1_n1015, position1_n1014, 
      position1_n1013, position1_n1012, position1_n1011, position1_n1010, 
      position1_n1009, position1_n1008, position1_n1007, position1_n1006, 
      position1_n1005, position1_n1004, position1_n1003, position1_n1002, 
      position1_n1001, position1_n1000, position1_n999, position1_n998, 
      position1_n997, position1_n996, position1_n995, position1_n994, 
      position1_n993, position1_n992, position1_n991, position1_n990, 
      position1_n989, position1_n988, position1_n987, position1_n986, 
      position1_n985, position1_n984, position1_n983, position1_n982, 
      position1_n981, position1_n980, position1_n979, position1_n978, 
      position1_n977, position1_n976, position1_n975, position1_n974, 
      position1_n973, position1_n972, position1_n971, position1_n970, 
      position1_n969, position1_n968, position1_n967, position1_n966, 
      position1_n965, position1_n964, position1_n963, position1_n962, 
      position1_n961, position1_n960, position1_n959, position1_n958, 
      position1_n957, position1_n956, position1_n955, position1_n954, 
      position1_n953, position1_n952, position1_n951, position1_n950, 
      position1_n949, position1_n948, position1_n947, position1_n946, 
      position1_n945, position1_n944, position1_n943, position1_n942, 
      position1_n941, position1_n940, position1_n939, position1_n938, 
      position1_n937, position1_n936, position1_n935, position1_n934, 
      position1_n933, position1_n932, position1_n931, position1_n930, 
      position1_n929, position1_n928, position1_n927, position1_n926, 
      position1_n925, position1_n924, position1_n923, position1_n922, 
      position1_n921, position1_n920, position1_n919, position1_n918, 
      position1_n917, position1_n916, position1_n915, position1_n914, 
      position1_n913, position1_n912, position1_n911, position1_n910, 
      position1_n909, position1_n908, position1_n907, position1_n906, 
      position1_n905, position1_n904, position1_n903, position1_n902, 
      position1_n901, position1_n900, position1_n899, position1_n898, 
      position1_n897, position1_n896, position1_n895, position1_n894, 
      position1_n893, position1_n892, position1_n891, position1_n890, 
      position1_n889, position1_n888, position1_n887, position1_n886, 
      position1_n885, position1_n884, position1_n883, position1_n882, 
      position1_n881, position1_n880, position1_n879, position1_n878, 
      position1_n877, position1_n876, position1_n875, position1_n874, 
      position1_n873, position1_n872, position1_n871, position1_n870, 
      position1_n869, position1_n868, position1_n867, position1_n866, 
      position1_n865, position1_n864, position1_n863, position1_n862, 
      position1_n861, position1_n860, position1_n859, position1_n858, 
      position1_n857, position1_n856, position1_n855, position1_n854, 
      position1_n853, position1_n852, position1_n851, position1_n850, 
      position1_n849, position1_n848, position1_n847, position1_n846, 
      position1_n845, position1_n844, position1_n843, position1_n842, 
      position1_n841, position1_n840, position1_n839, position1_n838, 
      position1_n837, position1_n836, position1_n835, position1_n834, 
      position1_n833, position1_n802, position1_n370, position1_n369, 
      position1_n368, position1_n367, position1_n366, position1_n365, 
      position1_n364, position1_n363, position1_n362, position1_n360, 
      position1_n358, position1_n357, position1_n356, position1_n353, 
      position1_n352, position1_n351, position1_n350, position1_n349, 
      position1_n348, position1_n347, position1_n346, position1_n344, 
      position1_n283, position1_dp_cluster_7_N314, position1_dp_cluster_6_N389,
      position1_N2460, position1_N2459, position1_N2458, position1_N2457, 
      position1_N2456, position1_N2455, position1_N2454, position1_N2453, 
      position1_N2452, position1_N2451, position1_N2450, position1_N2449, 
      position1_N2448, position1_N2447, position1_N2446, position1_N2445, 
      position1_N2413, position1_N2412, position1_N2411, position1_N2410, 
      position1_N2409, position1_N2408, position1_N2407, position1_N2406, 
      position1_N2405, position1_N2402, position1_N2401, position1_N2400, 
      position1_N2399, position1_N2398, position1_N2397, position1_N2396, 
      position1_N2395, position1_N2394, position1_N2391, position1_N2390, 
      position1_N2389, position1_N2388, position1_N2387, position1_N2386, 
      position1_N2385, position1_N2384, position1_N2383, position1_N2381, 
      position1_N2380, position1_N2379, position1_N2378, position1_N2377, 
      position1_N2376, position1_N2375, position1_N2374, position1_N2373, 
      position1_N2371, position1_N2370, position1_N2369, position1_N2368, 
      position1_N2367, position1_N2366, position1_N2365, position1_N2364, 
      position1_N2363, position1_N2362, position1_N2361, position1_N2360, 
      position1_N2359, position1_N2358, position1_N2357, position1_N2356, 
      position1_N2355, position1_N2354, position1_N2353, position1_N2352, 
      position1_N2326, position1_N2325, position1_N2324, position1_N2323, 
      position1_N2322, position1_N2321, position1_N2320, position1_N2319, 
      position1_N2318, position1_N2317, position1_N2316, position1_N2315, 
      position1_N2314, position1_N2313, position1_N2312, position1_N2311, 
      position1_N2310, position1_N2309, position1_N2308, position1_N2307, 
      position1_N2306, position1_N2305, position1_N2304, position1_N2303, 
      position1_N2300, position1_N2274, position1_N2273, position1_N2272, 
      position1_N2271, position1_N2270, position1_N2269, position1_N2268, 
      position1_N2267, position1_N2266, position1_N2265, position1_N2264, 
      position1_N2263, position1_N2262, position1_N2261, position1_N2260, 
      position1_N2259, position1_N2258, position1_N2257, position1_N2256, 
      position1_N2255, position1_N2254, position1_N2253, position1_N2252, 
      position1_N2248, position1_N2222, position1_N2221, position1_N2220, 
      position1_N2219, position1_N2218, position1_N2217, position1_N2216, 
      position1_N2215, position1_N2214, position1_N2213, position1_N2212, 
      position1_N2211, position1_N2210, position1_N2209, position1_N2208, 
      position1_N2207, position1_N2206, position1_N2205, position1_N2204, 
      position1_N2203, position1_N2202, position1_N2201, position1_N2196, 
      position1_N2170, position1_N2169, position1_N2168, position1_N2167, 
      position1_N2166, position1_N2165, position1_N2164, position1_N2163, 
      position1_N2162, position1_N2161, position1_N2160, position1_N2159, 
      position1_N2158, position1_N2157, position1_N2156, position1_N2155, 
      position1_N2154, position1_N2153, position1_N2152, position1_N2151, 
      position1_N2150, position1_N2144, position1_N2118, position1_N2117, 
      position1_N2116, position1_N2115, position1_N2114, position1_N2113, 
      position1_N2112, position1_N2111, position1_N2110, position1_N2109, 
      position1_N2108, position1_N2107, position1_N2106, position1_N2105, 
      position1_N2104, position1_N2103, position1_N2102, position1_N2101, 
      position1_N2100, position1_N2099, position1_N2094, position1_N2092, 
      position1_N2091, position1_N2090, position1_N2089, position1_N2088, 
      position1_N2087, position1_N2086, position1_N2085, position1_N2084, 
      position1_N2083, position1_N2082, position1_N2081, position1_N2080, 
      position1_N2079, position1_N2078, position1_N2077, position1_N2076, 
      position1_N2075, position1_N2074, position1_N2073, position1_N2072, 
      position1_N2071, position1_N2070, position1_N2069, position1_N2068, 
      position1_N2065, position1_N2064, position1_N2063, position1_N2062, 
      position1_N2061, position1_N2060, position1_N2059, position1_N2058, 
      position1_N2057, position1_N2056, position1_N2055, position1_N2054, 
      position1_N2053, position1_N2052, position1_N2051, position1_N2050, 
      position1_N2049, position1_N2040, position1_N2014, position1_N2013, 
      position1_N2012, position1_N2011, position1_N2010, position1_N2009, 
      position1_N2008, position1_N2007, position1_N2006, position1_N2005, 
      position1_N2004, position1_N2003, position1_N2002, position1_N2001, 
      position1_N2000, position1_N1999, position1_N1998, position1_N1997, 
      position1_N1990, position1_N1988, position1_N1987, position1_N1986, 
      position1_N1985, position1_N1984, position1_N1983, position1_N1982, 
      position1_N1981, position1_N1980, position1_N1979, position1_N1978, 
      position1_N1977, position1_N1976, position1_N1975, position1_N1974, 
      position1_N1973, position1_N1972, position1_N1971, position1_N1970, 
      position1_N1969, position1_N1968, position1_N1967, position1_N1966, 
      position1_N1965, position1_N1964, position1_N1962, position1_N1961, 
      position1_N1960, position1_N1959, position1_N1958, position1_N1957, 
      position1_N1956, position1_N1955, position1_N1954, position1_N1953, 
      position1_N1952, position1_N1951, position1_N1950, position1_N1949, 
      position1_N1948, position1_N1947, position1_N1946, position1_N1938, 
      position1_N1936, position1_N1935, position1_N1909, position1_N1908, 
      position1_N1907, position1_N1906, position1_N1905, position1_N1904, 
      position1_N1903, position1_N1902, position1_N1901, position1_N1900, 
      position1_N1899, position1_N1898, position1_N1897, position1_N1896, 
      position1_N1895, position1_N1894, position1_N1893, position1_N1892, 
      position1_N1891, position1_N1890, position1_N1889, position1_N1888, 
      position1_N1887, position1_N1886, position1_N1883, position1_N1857, 
      position1_N1856, position1_N1855, position1_N1854, position1_N1853, 
      position1_N1852, position1_N1851, position1_N1850, position1_N1849, 
      position1_N1848, position1_N1847, position1_N1846, position1_N1845, 
      position1_N1844, position1_N1843, position1_N1842, position1_N1841, 
      position1_N1840, position1_N1839, position1_N1838, position1_N1837, 
      position1_N1836, position1_N1835, position1_N1831, position1_N1805, 
      position1_N1804, position1_N1803, position1_N1802, position1_N1801, 
      position1_N1800, position1_N1799, position1_N1798, position1_N1797, 
      position1_N1796, position1_N1795, position1_N1794, position1_N1793, 
      position1_N1792, position1_N1791, position1_N1790, position1_N1789, 
      position1_N1788, position1_N1787, position1_N1786, position1_N1785, 
      position1_N1784, position1_N1779, position1_N1753, position1_N1752, 
      position1_N1751, position1_N1750, position1_N1749, position1_N1748, 
      position1_N1747, position1_N1746, position1_N1745, position1_N1744, 
      position1_N1743, position1_N1742, position1_N1741, position1_N1740, 
      position1_N1739, position1_N1738, position1_N1737, position1_N1736, 
      position1_N1735, position1_N1734, position1_N1733, position1_N1727, 
      position1_N1701, position1_N1700, position1_N1699, position1_N1698, 
      position1_N1697, position1_N1696, position1_N1695, position1_N1694, 
      position1_N1693, position1_N1692, position1_N1691, position1_N1690, 
      position1_N1689, position1_N1688, position1_N1687, position1_N1686, 
      position1_N1685, position1_N1684, position1_N1683, position1_N1682, 
      position1_N1677, position1_N1675, position1_N1674, position1_N1673, 
      position1_N1672, position1_N1671, position1_N1670, position1_N1669, 
      position1_N1668, position1_N1667, position1_N1666, position1_N1665, 
      position1_N1664, position1_N1663, position1_N1662, position1_N1661, 
      position1_N1660, position1_N1659, position1_N1658, position1_N1657, 
      position1_N1656, position1_N1655, position1_N1654, position1_N1653, 
      position1_N1652, position1_N1651, position1_N1648, position1_N1647, 
      position1_N1646, position1_N1645, position1_N1644, position1_N1643, 
      position1_N1642, position1_N1641, position1_N1640, position1_N1639, 
      position1_N1638, position1_N1637, position1_N1636, position1_N1635_port, 
      position1_N1634_port, position1_N1633_port, position1_N1632_port, 
      position1_N1623_port, position1_N1597_port, position1_N1596_port, 
      position1_N1595_port, position1_N1594_port, position1_N1593_port, 
      position1_N1592_port, position1_N1591_port, position1_N1590_port, 
      position1_N1589_port, position1_N1588_port, position1_N1587_port, 
      position1_N1586_port, position1_N1585_port, position1_N1584_port, 
      position1_N1583_port, position1_N1582_port, position1_N1581_port, 
      position1_N1580_port, position1_N1573_port, position1_N1571_port, 
      position1_N1570_port, position1_N1569_port, position1_N1568_port, 
      position1_N1567_port, position1_N1566_port, position1_N1565_port, 
      position1_N1564_port, position1_N1563_port, position1_N1562_port, 
      position1_N1561_port, position1_N1560_port, position1_N1559_port, 
      position1_N1558_port, position1_N1557_port, position1_N1556_port, 
      position1_N1555_port, position1_N1554_port, position1_N1553_port, 
      position1_N1552_port, position1_N1551_port, position1_N1550_port, 
      position1_N1549_port, position1_N1548_port, position1_N1547_port, 
      position1_N1545_port, position1_N1544_port, position1_N1543_port, 
      position1_N1542_port, position1_N1541_port, position1_N1540_port, 
      position1_N1539_port, position1_N1538_port, position1_N1537_port, 
      position1_N1536_port, position1_N1535_port, position1_N1534_port, 
      position1_N1533_port, position1_N1532_port, position1_N1531_port, 
      position1_N1530_port, position1_N1529_port, position1_N1521_port, 
      position1_N1519_port, position1_N1226_port, position1_N1225_port, 
      position1_N1224_port, position1_N1223_port, position1_N1222_port, 
      position1_N1221_port, position1_N1220_port, position1_N1219_port, 
      position1_N1218_port, position1_N1217_port, position1_N1216_port, 
      position1_N1215_port, position1_N1214_port, position1_N1213_port, 
      position1_N1212_port, position1_N1211_port, position1_N1210_port, 
      position1_N1209_port, position1_N1208_port, position1_N1207_port, 
      position1_N1206_port, position1_N1205_port, position1_N1204_port, 
      position1_N1203_port, position1_N1202_port, position1_N1201_port, 
      position1_N1200_port, position1_N1199_port, position1_N1198_port, 
      position1_N1197_port, position1_N1196_port, position1_N1195_port, 
      position1_N1194_port, position1_N1193_port, position1_N1192_port, 
      position1_N1191_port, position1_N1190_port, position1_N1189_port, 
      position1_N1188_port, position1_N1187_port, position1_N1186_port, 
      position1_N1185_port, position1_N1184_port, position1_N1183_port, 
      position1_N1182_port, position1_N1181_port, position1_N1180_port, 
      position1_N1179_port, position1_N1178_port, position1_N1177_port, 
      position1_N1003_port, position1_N1002_port, position1_N1001_port, 
      position1_N1000_port, position1_N999_port, position1_N998_port, 
      position1_N997_port, position1_N996_port, position1_N995_port, 
      position1_N994_port, position1_N993_port, position1_N992_port, 
      position1_N991_port, position1_N990_port, position1_N989_port, 
      position1_N988_port, position1_N987_port, position1_N986_port, 
      position1_N985_port, position1_N984_port, position1_N983_port, 
      position1_N982_port, position1_N981_port, position1_N980_port, 
      position1_N928_port, position1_N927_port, position1_N926_port, 
      position1_N925_port, position1_N924_port, position1_N923_port, 
      position1_N922_port, position1_N921_port, position1_N920_port, 
      position1_N919_port, position1_N918_port, position1_N917_port, 
      position1_N916_port, position1_N915_port, position1_N914_port, 
      position1_N913_port, position1_N912_port, position1_N911_port, 
      position1_N910_port, position1_N909_port, position1_N908_port, 
      position1_N907_port, position1_N906_port, position1_N905_port, 
      position1_N656, position1_N655, position1_N654, position1_N653, 
      position1_N652, position1_N651, position1_N650, position1_N649, 
      position1_N648, position1_N647, position1_N646, position1_N645, 
      position1_N644, position1_N643, position1_N642, position1_N641, 
      position1_N640, position1_N639, position1_N638, position1_N637, 
      position1_N636, position1_N635, position1_N634, position1_N633, 
      position1_N632, position1_N631, position1_N630, position1_N629, 
      position1_N628, position1_N627, position1_N626, position1_N625, 
      position1_N624, position1_N623, position1_N622, position1_N621, 
      position1_N620, position1_N619, position1_N618, position1_N617, 
      position1_N616, position1_N615, position1_N614, position1_N613, 
      position1_N612, position1_N611, position1_N610, position1_N609, 
      position1_N608, position1_N607, position1_N606, position1_N605, 
      position1_N604, position1_N603, position1_N602, position1_N601, 
      position1_N600, position1_N599, position1_N598, position1_N597, 
      position1_N596, position1_N595, position1_N594, position1_N593, 
      position1_N592, position1_N591, position1_N590, position1_N577, 
      position1_N576, position1_N575, position1_N574, position1_N573, 
      position1_N572, position1_N571, position1_N570, position1_N569, 
      position1_N568, position1_N567, position1_N566, position1_N565, 
      position1_N564, position1_N563, position1_N562, position1_N560, 
      position1_N559, position1_N558, position1_N557, position1_N556, 
      position1_N555, position1_N554, position1_N553, position1_N552, 
      position1_N551, position1_N550, position1_N549, position1_N548, 
      position1_N547, position1_N546, position1_N545, position1_N544, 
      position1_N543, position1_N542, position1_N541, position1_N540, 
      position1_N539, position1_N538, position1_N537, position1_N536, 
      position1_N535, position1_N509, position1_N508, position1_N507, 
      position1_N506, position1_N505, position1_N504, position1_N503, 
      position1_N502, position1_N501, position1_N500, position1_N499, 
      position1_N498, position1_N497, position1_N496, position1_N495, 
      position1_N494, position1_N493, position1_N492, position1_N491, 
      position1_N490, position1_N489, position1_N488, position1_N487, 
      position1_N486, position1_N485, position1_N447, position1_N446, 
      position1_N445, position1_N444, position1_N443, position1_N442, 
      position1_N441, position1_N440, position1_N439, position1_N438, 
      position1_N437, position1_N436, position1_N435, position1_N434, 
      position1_N433, position1_N432, position1_N431, position1_N429, 
      position1_N428, position1_N427, position1_N426, position1_N425, 
      position1_N424, position1_N423, position1_N422, position1_N421, 
      position1_N420, position1_N419, position1_N418, position1_N417, 
      position1_N416, position1_N415, position1_N414, position1_N413, 
      position1_N412, position1_N411, position1_N410, position1_N409, 
      position1_N408, position1_N407, position1_N406, position1_N379, 
      position1_N378, position1_N377, position1_N376, position1_N375, 
      position1_N374, position1_N373, position1_N372, position1_N371, 
      position1_N370_port, position1_N369_port, position1_N368_port, 
      position1_N367_port, position1_N366_port, position1_N365_port, 
      position1_N364_port, position1_N363_port, position1_N362_port, 
      position1_N361, position1_N360_port, position1_N359, position1_N358_port,
      position1_N357_port, position1_N356_port, position1_N355, position1_N354,
      position1_N353_port, position1_N352_port, position1_N351_port, 
      position1_N350_port, position1_N349_port, position1_N348_port, 
      position1_N347_port, position1_N346_port, position1_N345, 
      position1_N344_port, position1_N343, position1_N342, position1_N341, 
      position1_N340, position1_N339, position1_N338, position1_N337, 
      position1_N336, position1_N335, position1_N334, position1_N333, 
      position1_N332, position1_N331, position1_N304, position1_N303, 
      position1_N302, position1_N301, position1_N300, position1_N299, 
      position1_N298, position1_N297, position1_N296, position1_N295, 
      position1_N294, position1_N293, position1_N292, position1_N291, 
      position1_N290, position1_N289, position1_N288, position1_N287, 
      position1_N286, position1_N285, position1_N284, position1_N283_port, 
      position1_N282, position1_N281, position1_N280, position1_N267, 
      position1_N224, position1_N223, position1_N222, position1_N221, 
      position1_N220, position1_N219, position1_N218, position1_N217, 
      position1_N216, position1_N215, position1_N214, position1_N213, 
      position1_N212, position1_N211, position1_N210, position1_N209, 
      position1_N208, position1_N207, position1_N206, position1_quot_y_0_port, 
      position1_quot_y_1_port, position1_quot_y_2_port, position1_quot_y_3_port
      , position1_quot_y_4_port, position1_quot_y_5_port, 
      position1_quot_y_6_port, position1_quot_y_7_port, position1_quot_y_8_port
      , position1_quot_x_0_port, position1_quot_x_1_port, 
      position1_quot_x_2_port, position1_quot_x_3_port, position1_quot_x_4_port
      , position1_quot_x_5_port, position1_quot_x_6_port, 
      position1_quot_x_7_port, position1_quot_x_8_port, position1_N194, 
      position1_N193, position1_N104, position1_N103, position1_N102, 
      position1_N101, position1_N100, position1_N99, position1_N98, 
      position1_N97, position1_N95, position1_N94, position1_N93, position1_N91
      , position1_N89, position1_N88, position1_N87, position1_N86, 
      position1_N85, position1_N84, position1_N83, position1_N82, position1_N81
      , position1_state_0_port, position1_state_1_port, 
      position1_count_img_0_port, position1_count_img_1_port, 
      position1_count_img_2_port, position1_count_img_3_port, 
      position1_count_img_4_port, position1_count_img_5_port, 
      position1_count_img_6_port, position1_count_img_7_port, 
      position1_count_img_8_port, position1_count_img_9_port, 
      position1_count_img_10_port, position1_count_img_11_port, 
      position1_count_img_12_port, position1_count_img_13_port, 
      position1_count_img_14_port, position1_count_img_15_port, 
      position1_count_img_16_port, position1_count_img_17_port, 
      position1_count_img_18_port, position1_count_img_19_port, 
      position1_y_sum_1_port, position1_y_sum_2_port, position1_y_sum_3_port, 
      position1_y_sum_4_port, position1_y_sum_5_port, position1_y_sum_6_port, 
      position1_y_sum_7_port, position1_y_sum_8_port, position1_y_sum_9_port, 
      position1_y_sum_10_port, position1_y_sum_11_port, position1_y_sum_12_port
      , position1_y_sum_13_port, position1_y_sum_14_port, 
      position1_y_sum_15_port, position1_y_sum_16_port, position1_y_sum_17_port
      , position1_y_sum_18_port, position1_y_sum_19_port, 
      position1_y_sum_20_port, position1_y_sum_21_port, position1_y_sum_22_port
      , position1_y_sum_23_port, position1_y_sum_24_port, 
      position1_x_sum_1_port, position1_x_sum_2_port, position1_x_sum_3_port, 
      position1_x_sum_4_port, position1_x_sum_5_port, position1_x_sum_6_port, 
      position1_x_sum_7_port, position1_x_sum_8_port, position1_x_sum_9_port, 
      position1_x_sum_10_port, position1_x_sum_11_port, position1_x_sum_12_port
      , position1_x_sum_13_port, position1_x_sum_14_port, 
      position1_x_sum_15_port, position1_x_sum_16_port, position1_x_sum_17_port
      , position1_x_sum_18_port, position1_x_sum_19_port, 
      position1_x_sum_20_port, position1_x_sum_21_port, position1_x_sum_22_port
      , position1_x_sum_23_port, position1_x_sum_24_port, position1_gi_0_port, 
      position1_gi_1_port, position1_gi_2_port, position1_gi_3_port, 
      position1_gi_4_port, position1_gi_5_port, position1_gi_6_port, 
      position1_gi_7_port, position1_r406_carry_1_port, 
      position1_r406_carry_2_port, position1_r406_carry_3_port, 
      position1_r406_carry_4_port, position1_r406_carry_5_port, 
      position1_r406_carry_6_port, position1_r406_carry_7_port, 
      position1_r406_carry_8_port, position1_r406_carry_9_port, 
      position1_r406_carry_10_port, position1_r406_carry_11_port, 
      position1_r406_carry_12_port, position1_r406_carry_13_port, 
      position1_r406_carry_14_port, position1_r406_carry_15_port, 
      position1_r406_carry_16_port, position1_r406_carry_17_port, 
      position1_r406_carry_18_port, position1_r406_carry_19_port, 
      position1_r406_carry_20_port, position1_r406_carry_21_port, 
      position1_r406_carry_22_port, position1_r406_carry_23_port, 
      position1_r406_carry_24_port, position1_r409_carry_1_port, 
      position1_r409_carry_2_port, position1_r409_carry_3_port, 
      position1_r409_carry_4_port, position1_r409_carry_5_port, 
      position1_r409_carry_6_port, position1_r409_carry_7_port, 
      position1_r409_carry_8_port, position1_r409_carry_9_port, 
      position1_r409_carry_10_port, position1_r409_carry_11_port, 
      position1_r409_carry_12_port, position1_r409_carry_13_port, 
      position1_r409_carry_14_port, position1_r409_carry_15_port, 
      position1_r409_carry_16_port, position1_r409_carry_17_port, 
      position1_r409_carry_18_port, position1_r409_carry_19_port, 
      position1_r409_carry_20_port, position1_r409_carry_21_port, 
      position1_r409_carry_22_port, position1_r409_carry_23_port, 
      position1_r409_carry_24_port, position1_r412_carry_1_port, 
      position1_r412_carry_2_port, position1_r412_carry_3_port, 
      position1_r412_carry_4_port, position1_r412_carry_5_port, 
      position1_r412_carry_6_port, position1_r412_carry_7_port, 
      position1_r412_carry_8_port, position1_r412_carry_9_port, 
      position1_r412_carry_10_port, position1_r412_carry_11_port, 
      position1_r412_carry_12_port, position1_r412_carry_13_port, 
      position1_r412_carry_14_port, position1_r412_carry_15_port, 
      position1_r412_carry_16_port, position1_r412_carry_17_port, 
      position1_r412_carry_18_port, position1_r412_carry_19_port, 
      position1_r412_carry_20_port, position1_r412_carry_21_port, 
      position1_r412_carry_22_port, position1_r412_carry_23_port, 
      position1_r412_carry_24_port, position1_r413_carry_1_port, 
      position1_r413_carry_2_port, position1_r413_carry_3_port, 
      position1_r413_carry_4_port, position1_r413_carry_5_port, 
      position1_r413_carry_6_port, position1_r413_carry_7_port, 
      position1_r413_carry_8_port, position1_r413_carry_9_port, 
      position1_r413_carry_10_port, position1_r413_carry_11_port, 
      position1_r413_carry_12_port, position1_r413_carry_13_port, 
      position1_r413_carry_14_port, position1_r413_carry_15_port, 
      position1_r413_carry_16_port, position1_r413_carry_17_port, 
      position1_r413_carry_18_port, position1_r413_carry_19_port, 
      position1_r413_carry_20_port, position1_r413_carry_21_port, 
      position1_r413_carry_22_port, position1_r413_carry_23_port, 
      position1_r413_carry_24_port, position1_r416_carry_2_port, 
      position1_r416_carry_3_port, position1_r416_carry_4_port, 
      position1_r416_carry_5_port, position1_r416_carry_6_port, 
      position1_r416_carry_7_port, position1_r416_carry_8_port, 
      position1_r416_carry_9_port, position1_r416_carry_10_port, 
      position1_r416_carry_11_port, position1_r416_carry_12_port, 
      position1_r416_carry_13_port, position1_r416_carry_14_port, 
      position1_r416_carry_15_port, position1_r416_carry_16_port, 
      position1_r416_carry_17_port, position1_r457_carry_2_port, 
      position1_r457_carry_3_port, position1_r457_carry_4_port, 
      position1_r457_carry_5_port, position1_r457_carry_6_port, 
      position1_r457_carry_7_port, position1_r457_carry_8_port, 
      position1_r457_carry_9_port, position1_r457_carry_10_port, 
      position1_r457_carry_11_port, position1_r457_carry_12_port, 
      position1_r457_carry_13_port, position1_r457_carry_14_port, 
      position1_r457_carry_15_port, position1_r457_carry_16_port, 
      position1_r457_carry_17_port, position1_r458_carry_3_port, 
      position1_r458_carry_4_port, position1_r458_carry_5_port, 
      position1_r458_carry_6_port, position1_r458_carry_7_port, 
      position1_r458_carry_8_port, position1_r458_carry_9_port, 
      position1_r458_carry_10_port, position1_r458_carry_11_port, 
      position1_r458_carry_12_port, position1_r458_carry_13_port, 
      position1_r458_carry_14_port, position1_r458_carry_15_port, 
      position1_r458_carry_16_port, position1_r458_carry_17_port, 
      position1_add_161_carry_2_port, position1_add_161_carry_3_port, 
      position1_add_161_carry_4_port, position1_add_161_carry_5_port, 
      position1_add_161_carry_6_port, position1_add_161_carry_7_port, 
      position1_add_161_carry_8_port, position1_add_161_carry_9_port, 
      position1_add_161_carry_10_port, position1_add_161_carry_11_port, 
      position1_add_161_carry_12_port, position1_add_161_carry_13_port, 
      position1_add_161_carry_14_port, position1_add_161_carry_15_port, 
      position1_add_161_carry_16_port, position1_add_161_carry_17_port, 
      position1_add_161_carry_18_port, position1_add_161_carry_19_port, 
      position1_sub_216_carry_9_port, position1_sub_216_carry_10_port, 
      position1_sub_216_carry_11_port, position1_sub_216_carry_12_port, 
      position1_sub_216_carry_13_port, position1_sub_216_carry_14_port, 
      position1_sub_216_carry_15_port, position1_sub_216_carry_16_port, 
      position1_sub_216_carry_17_port, position1_sub_216_carry_18_port, 
      position1_sub_216_carry_19_port, position1_sub_216_carry_20_port, 
      position1_sub_216_carry_21_port, position1_sub_216_carry_22_port, 
      position1_sub_216_carry_23_port, position1_sub_216_carry_24_port, 
      position1_sub_216_I2_carry_8_port, position1_sub_216_I2_carry_9_port, 
      position1_sub_216_I2_carry_10_port, position1_sub_216_I2_carry_11_port, 
      position1_sub_216_I2_carry_12_port, position1_sub_216_I2_carry_13_port, 
      position1_sub_216_I2_carry_14_port, position1_sub_216_I2_carry_15_port, 
      position1_sub_216_I2_carry_16_port, position1_sub_216_I2_carry_17_port, 
      position1_sub_216_I2_carry_18_port, position1_sub_216_I2_carry_19_port, 
      position1_sub_216_I2_carry_20_port, position1_sub_216_I2_carry_21_port, 
      position1_sub_216_I2_carry_22_port, position1_sub_216_I2_carry_23_port, 
      position1_sub_216_I2_carry_24_port, position1_sub_216_I3_carry_7_port, 
      position1_sub_216_I3_carry_8_port, position1_sub_216_I3_carry_9_port, 
      position1_sub_216_I3_carry_10_port, position1_sub_216_I3_carry_11_port, 
      position1_sub_216_I3_carry_12_port, position1_sub_216_I3_carry_13_port, 
      position1_sub_216_I3_carry_14_port, position1_sub_216_I3_carry_15_port, 
      position1_sub_216_I3_carry_16_port, position1_sub_216_I3_carry_17_port, 
      position1_sub_216_I3_carry_18_port, position1_sub_216_I3_carry_19_port, 
      position1_sub_216_I3_carry_20_port, position1_sub_216_I3_carry_21_port, 
      position1_sub_216_I3_carry_22_port, position1_sub_216_I3_carry_23_port, 
      position1_sub_216_I3_carry_24_port, position1_sub_216_I4_carry_6_port, 
      position1_sub_216_I4_carry_7_port, position1_sub_216_I4_carry_8_port, 
      position1_sub_216_I4_carry_9_port, position1_sub_216_I4_carry_10_port, 
      position1_sub_216_I4_carry_11_port, position1_sub_216_I4_carry_12_port, 
      position1_sub_216_I4_carry_13_port, position1_sub_216_I4_carry_14_port, 
      position1_sub_216_I4_carry_15_port, position1_sub_216_I4_carry_16_port, 
      position1_sub_216_I4_carry_17_port, position1_sub_216_I4_carry_18_port, 
      position1_sub_216_I4_carry_19_port, position1_sub_216_I4_carry_20_port, 
      position1_sub_216_I4_carry_21_port, position1_sub_216_I4_carry_22_port, 
      position1_sub_216_I4_carry_23_port, position1_sub_216_I4_carry_24_port, 
      position1_sub_216_I5_carry_5_port, position1_sub_216_I5_carry_6_port, 
      position1_sub_216_I5_carry_7_port, position1_sub_216_I5_carry_8_port, 
      position1_sub_216_I5_carry_9_port, position1_sub_216_I5_carry_10_port, 
      position1_sub_216_I5_carry_11_port, position1_sub_216_I5_carry_12_port, 
      position1_sub_216_I5_carry_13_port, position1_sub_216_I5_carry_14_port, 
      position1_sub_216_I5_carry_15_port, position1_sub_216_I5_carry_16_port, 
      position1_sub_216_I5_carry_17_port, position1_sub_216_I5_carry_18_port, 
      position1_sub_216_I5_carry_19_port, position1_sub_216_I5_carry_20_port, 
      position1_sub_216_I5_carry_21_port, position1_sub_216_I5_carry_22_port, 
      position1_sub_216_I5_carry_23_port, position1_sub_216_I5_carry_24_port, 
      position1_sub_216_I6_carry_4_port, position1_sub_216_I6_carry_5_port, 
      position1_sub_216_I6_carry_6_port, position1_sub_216_I6_carry_7_port, 
      position1_sub_216_I6_carry_8_port, position1_sub_216_I6_carry_9_port, 
      position1_sub_216_I6_carry_10_port, position1_sub_216_I6_carry_11_port, 
      position1_sub_216_I6_carry_12_port, position1_sub_216_I6_carry_13_port, 
      position1_sub_216_I6_carry_14_port, position1_sub_216_I6_carry_15_port, 
      position1_sub_216_I6_carry_16_port, position1_sub_216_I6_carry_17_port, 
      position1_sub_216_I6_carry_18_port, position1_sub_216_I6_carry_19_port, 
      position1_sub_216_I6_carry_20_port, position1_sub_216_I6_carry_21_port, 
      position1_sub_216_I6_carry_22_port, position1_sub_216_I6_carry_23_port, 
      position1_sub_216_I6_carry_24_port, position1_sub_216_I7_carry_3_port, 
      position1_sub_216_I7_carry_4_port, position1_sub_216_I7_carry_5_port, 
      position1_sub_216_I7_carry_6_port, position1_sub_216_I7_carry_7_port, 
      position1_sub_216_I7_carry_8_port, position1_sub_216_I7_carry_9_port, 
      position1_sub_216_I7_carry_10_port, position1_sub_216_I7_carry_11_port, 
      position1_sub_216_I7_carry_12_port, position1_sub_216_I7_carry_13_port, 
      position1_sub_216_I7_carry_14_port, position1_sub_216_I7_carry_15_port, 
      position1_sub_216_I7_carry_16_port, position1_sub_216_I7_carry_17_port, 
      position1_sub_216_I7_carry_18_port, position1_sub_216_I7_carry_19_port, 
      position1_sub_216_I7_carry_20_port, position1_sub_216_I7_carry_21_port, 
      position1_sub_216_I7_carry_22_port, position1_sub_216_I7_carry_23_port, 
      position1_sub_216_I7_carry_24_port, position1_sub_216_I8_carry_2_port, 
      position1_sub_216_I8_carry_3_port, position1_sub_216_I8_carry_4_port, 
      position1_sub_216_I8_carry_5_port, position1_sub_216_I8_carry_6_port, 
      position1_sub_216_I8_carry_7_port, position1_sub_216_I8_carry_8_port, 
      position1_sub_216_I8_carry_9_port, position1_sub_216_I8_carry_10_port, 
      position1_sub_216_I8_carry_11_port, position1_sub_216_I8_carry_12_port, 
      position1_sub_216_I8_carry_13_port, position1_sub_216_I8_carry_14_port, 
      position1_sub_216_I8_carry_15_port, position1_sub_216_I8_carry_16_port, 
      position1_sub_216_I8_carry_17_port, position1_sub_216_I8_carry_18_port, 
      position1_sub_216_I8_carry_19_port, position1_sub_216_I8_carry_20_port, 
      position1_sub_216_I8_carry_21_port, position1_sub_216_I8_carry_22_port, 
      position1_sub_216_I8_carry_23_port, position1_sub_226_carry_9_port, 
      position1_sub_226_carry_10_port, position1_sub_226_carry_11_port, 
      position1_sub_226_carry_12_port, position1_sub_226_carry_13_port, 
      position1_sub_226_carry_14_port, position1_sub_226_carry_15_port, 
      position1_sub_226_carry_16_port, position1_sub_226_carry_17_port, 
      position1_sub_226_carry_18_port, position1_sub_226_carry_19_port, 
      position1_sub_226_carry_20_port, position1_sub_226_carry_21_port, 
      position1_sub_226_carry_22_port, position1_sub_226_carry_23_port, 
      position1_sub_226_carry_24_port, position1_sub_226_I2_carry_8_port, 
      position1_sub_226_I2_carry_9_port, position1_sub_226_I2_carry_10_port, 
      position1_sub_226_I2_carry_11_port, position1_sub_226_I2_carry_12_port, 
      position1_sub_226_I2_carry_13_port, position1_sub_226_I2_carry_14_port, 
      position1_sub_226_I2_carry_15_port, position1_sub_226_I2_carry_16_port, 
      position1_sub_226_I2_carry_17_port, position1_sub_226_I2_carry_18_port, 
      position1_sub_226_I2_carry_19_port, position1_sub_226_I2_carry_20_port, 
      position1_sub_226_I2_carry_21_port, position1_sub_226_I2_carry_22_port, 
      position1_sub_226_I2_carry_23_port, position1_sub_226_I2_carry_24_port, 
      position1_sub_226_I3_carry_7_port, position1_sub_226_I3_carry_8_port, 
      position1_sub_226_I3_carry_9_port, position1_sub_226_I3_carry_10_port, 
      position1_sub_226_I3_carry_11_port, position1_sub_226_I3_carry_12_port, 
      position1_sub_226_I3_carry_13_port, position1_sub_226_I3_carry_14_port, 
      position1_sub_226_I3_carry_15_port, position1_sub_226_I3_carry_16_port, 
      position1_sub_226_I3_carry_17_port, position1_sub_226_I3_carry_18_port, 
      position1_sub_226_I3_carry_19_port, position1_sub_226_I3_carry_20_port, 
      position1_sub_226_I3_carry_21_port, position1_sub_226_I3_carry_22_port, 
      position1_sub_226_I3_carry_23_port, position1_sub_226_I3_carry_24_port, 
      position1_sub_226_I4_carry_6_port, position1_sub_226_I4_carry_7_port, 
      position1_sub_226_I4_carry_8_port, position1_sub_226_I4_carry_9_port, 
      position1_sub_226_I4_carry_10_port, position1_sub_226_I4_carry_11_port, 
      position1_sub_226_I4_carry_12_port, position1_sub_226_I4_carry_13_port, 
      position1_sub_226_I4_carry_14_port, position1_sub_226_I4_carry_15_port, 
      position1_sub_226_I4_carry_16_port, position1_sub_226_I4_carry_17_port, 
      position1_sub_226_I4_carry_18_port, position1_sub_226_I4_carry_19_port, 
      position1_sub_226_I4_carry_20_port, position1_sub_226_I4_carry_21_port, 
      position1_sub_226_I4_carry_22_port, position1_sub_226_I4_carry_23_port, 
      position1_sub_226_I4_carry_24_port, position1_sub_226_I5_carry_5_port, 
      position1_sub_226_I5_carry_6_port, position1_sub_226_I5_carry_7_port, 
      position1_sub_226_I5_carry_8_port, position1_sub_226_I5_carry_9_port, 
      position1_sub_226_I5_carry_10_port, position1_sub_226_I5_carry_11_port, 
      position1_sub_226_I5_carry_12_port, position1_sub_226_I5_carry_13_port, 
      position1_sub_226_I5_carry_14_port, position1_sub_226_I5_carry_15_port, 
      position1_sub_226_I5_carry_16_port, position1_sub_226_I5_carry_17_port, 
      position1_sub_226_I5_carry_18_port, position1_sub_226_I5_carry_19_port, 
      position1_sub_226_I5_carry_20_port, position1_sub_226_I5_carry_21_port, 
      position1_sub_226_I5_carry_22_port, position1_sub_226_I5_carry_23_port, 
      position1_sub_226_I5_carry_24_port, position1_sub_226_I6_carry_4_port, 
      position1_sub_226_I6_carry_5_port, position1_sub_226_I6_carry_6_port, 
      position1_sub_226_I6_carry_7_port, position1_sub_226_I6_carry_8_port, 
      position1_sub_226_I6_carry_9_port, position1_sub_226_I6_carry_10_port, 
      position1_sub_226_I6_carry_11_port, position1_sub_226_I6_carry_12_port, 
      position1_sub_226_I6_carry_13_port, position1_sub_226_I6_carry_14_port, 
      position1_sub_226_I6_carry_15_port, position1_sub_226_I6_carry_16_port, 
      position1_sub_226_I6_carry_17_port, position1_sub_226_I6_carry_18_port, 
      position1_sub_226_I6_carry_19_port, position1_sub_226_I6_carry_20_port, 
      position1_sub_226_I6_carry_21_port, position1_sub_226_I6_carry_22_port, 
      position1_sub_226_I6_carry_23_port, position1_sub_226_I6_carry_24_port, 
      position1_sub_226_I7_carry_3_port, position1_sub_226_I7_carry_4_port, 
      position1_sub_226_I7_carry_5_port, position1_sub_226_I7_carry_6_port, 
      position1_sub_226_I7_carry_7_port, position1_sub_226_I7_carry_8_port, 
      position1_sub_226_I7_carry_9_port, position1_sub_226_I7_carry_10_port, 
      position1_sub_226_I7_carry_11_port, position1_sub_226_I7_carry_12_port, 
      position1_sub_226_I7_carry_13_port, position1_sub_226_I7_carry_14_port, 
      position1_sub_226_I7_carry_15_port, position1_sub_226_I7_carry_16_port, 
      position1_sub_226_I7_carry_17_port, position1_sub_226_I7_carry_18_port, 
      position1_sub_226_I7_carry_19_port, position1_sub_226_I7_carry_20_port, 
      position1_sub_226_I7_carry_21_port, position1_sub_226_I7_carry_22_port, 
      position1_sub_226_I7_carry_23_port, position1_sub_226_I7_carry_24_port, 
      position1_sub_226_I8_carry_2_port, position1_sub_226_I8_carry_3_port, 
      position1_sub_226_I8_carry_4_port, position1_sub_226_I8_carry_5_port, 
      position1_sub_226_I8_carry_6_port, position1_sub_226_I8_carry_7_port, 
      position1_sub_226_I8_carry_8_port, position1_sub_226_I8_carry_9_port, 
      position1_sub_226_I8_carry_10_port, position1_sub_226_I8_carry_11_port, 
      position1_sub_226_I8_carry_12_port, position1_sub_226_I8_carry_13_port, 
      position1_sub_226_I8_carry_14_port, position1_sub_226_I8_carry_15_port, 
      position1_sub_226_I8_carry_16_port, position1_sub_226_I8_carry_17_port, 
      position1_sub_226_I8_carry_18_port, position1_sub_226_I8_carry_19_port, 
      position1_sub_226_I8_carry_20_port, position1_sub_226_I8_carry_21_port, 
      position1_sub_226_I8_carry_22_port, position1_sub_226_I8_carry_23_port, 
      position1_sub_250_carry_2_port, position1_sub_250_carry_3_port, 
      position1_sub_250_carry_4_port, position1_sub_250_carry_5_port, 
      position1_sub_250_carry_6_port, position1_sub_250_carry_7_port, 
      position1_sub_250_3_carry_2_port, position1_sub_250_3_carry_3_port, 
      position1_sub_250_3_carry_4_port, position1_sub_250_3_carry_5_port, 
      position1_sub_250_3_carry_6_port, position1_sub_250_3_carry_7_port, 
      position1_add_250_carry_2_port, position1_add_250_carry_3_port, 
      position1_add_250_carry_4_port, position1_add_250_carry_5_port, 
      position1_add_250_carry_6_port, position1_add_250_carry_7_port, 
      position1_add_250_carry_8_port, position1_add_250_2_carry_2_port, 
      position1_add_250_2_carry_3_port, position1_add_250_2_carry_4_port, 
      position1_add_250_2_carry_5_port, position1_add_250_2_carry_6_port, 
      position1_add_250_2_carry_7_port, position1_add_250_2_carry_8_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_0_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_1_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_2_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_3_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_4_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_5_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_6_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_7_port, 
      position1_dp_cluster_0_mult_add_196_aco_PROD_not_8_port, 
      position1_dp_cluster_0_add_196_aco_carry_1_port, 
      position1_dp_cluster_0_add_196_aco_carry_2_port, 
      position1_dp_cluster_0_add_196_aco_carry_3_port, 
      position1_dp_cluster_0_add_196_aco_carry_4_port, 
      position1_dp_cluster_0_add_196_aco_carry_5_port, 
      position1_dp_cluster_0_add_196_aco_carry_6_port, 
      position1_dp_cluster_0_add_196_aco_carry_7_port, 
      position1_dp_cluster_0_add_196_aco_carry_8_port, 
      position1_dp_cluster_0_add_196_aco_carry_9_port, 
      position1_dp_cluster_0_add_196_aco_carry_10_port, 
      position1_dp_cluster_0_add_196_aco_carry_11_port, 
      position1_dp_cluster_0_add_196_aco_carry_12_port, 
      position1_dp_cluster_0_add_196_aco_carry_13_port, 
      position1_dp_cluster_0_add_196_aco_carry_14_port, 
      position1_dp_cluster_0_add_196_aco_carry_15_port, 
      position1_dp_cluster_0_add_196_aco_carry_16_port, 
      position1_dp_cluster_0_add_196_aco_carry_17_port, 
      position1_dp_cluster_0_add_196_aco_carry_18_port, 
      position1_dp_cluster_0_add_196_aco_carry_19_port, 
      position1_dp_cluster_0_add_196_aco_carry_20_port, 
      position1_dp_cluster_0_add_196_aco_carry_21_port, 
      position1_dp_cluster_0_add_196_aco_carry_22_port, 
      position1_dp_cluster_0_add_196_aco_carry_23_port, 
      position1_dp_cluster_0_add_196_aco_carry_24_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_0_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_1_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_2_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_3_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_4_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_5_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_6_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_7_port, 
      position1_dp_cluster_1_mult_add_197_aco_PROD_not_8_port, 
      position1_dp_cluster_1_add_197_aco_carry_1_port, 
      position1_dp_cluster_1_add_197_aco_carry_2_port, 
      position1_dp_cluster_1_add_197_aco_carry_3_port, 
      position1_dp_cluster_1_add_197_aco_carry_4_port, 
      position1_dp_cluster_1_add_197_aco_carry_5_port, 
      position1_dp_cluster_1_add_197_aco_carry_6_port, 
      position1_dp_cluster_1_add_197_aco_carry_7_port, 
      position1_dp_cluster_1_add_197_aco_carry_8_port, 
      position1_dp_cluster_1_add_197_aco_carry_9_port, 
      position1_dp_cluster_1_add_197_aco_carry_10_port, 
      position1_dp_cluster_1_add_197_aco_carry_11_port, 
      position1_dp_cluster_1_add_197_aco_carry_12_port, 
      position1_dp_cluster_1_add_197_aco_carry_13_port, 
      position1_dp_cluster_1_add_197_aco_carry_14_port, 
      position1_dp_cluster_1_add_197_aco_carry_15_port, 
      position1_dp_cluster_1_add_197_aco_carry_16_port, 
      position1_dp_cluster_1_add_197_aco_carry_17_port, 
      position1_dp_cluster_1_add_197_aco_carry_18_port, 
      position1_dp_cluster_1_add_197_aco_carry_19_port, 
      position1_dp_cluster_1_add_197_aco_carry_20_port, 
      position1_dp_cluster_1_add_197_aco_carry_21_port, 
      position1_dp_cluster_1_add_197_aco_carry_22_port, 
      position1_dp_cluster_1_add_197_aco_carry_23_port, 
      position1_dp_cluster_1_add_197_aco_carry_24_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_2_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_3_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_4_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_5_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_6_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_7_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_8_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_9_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_10_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_11_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_12_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_13_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_14_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_15_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_16_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_17_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_18_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_19_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_20_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_21_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_22_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_23_port, 
      position1_dp_cluster_2_add_0_root_add_189_3_carry_24_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_2_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_3_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_4_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_5_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_6_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_7_port, 
      position1_dp_cluster_3_add_1_root_add_188_3_carry_8_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_2_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_3_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_4_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_5_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_6_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_7_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_8_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_9_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_10_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_11_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_12_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_13_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_14_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_15_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_16_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_17_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_18_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_19_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_20_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_21_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_22_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_23_port, 
      position1_dp_cluster_3_add_0_root_add_188_3_carry_24_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_0_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_1_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_2_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_3_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_4_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_5_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_6_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_7_port, 
      position1_dp_cluster_4_mult_add_178_aco_PROD_not_8_port, 
      position1_dp_cluster_4_add_178_aco_carry_1_port, 
      position1_dp_cluster_4_add_178_aco_carry_2_port, 
      position1_dp_cluster_4_add_178_aco_carry_3_port, 
      position1_dp_cluster_4_add_178_aco_carry_4_port, 
      position1_dp_cluster_4_add_178_aco_carry_5_port, 
      position1_dp_cluster_4_add_178_aco_carry_6_port, 
      position1_dp_cluster_4_add_178_aco_carry_7_port, 
      position1_dp_cluster_4_add_178_aco_carry_8_port, 
      position1_dp_cluster_4_add_178_aco_carry_9_port, 
      position1_dp_cluster_4_add_178_aco_carry_10_port, 
      position1_dp_cluster_4_add_178_aco_carry_11_port, 
      position1_dp_cluster_4_add_178_aco_carry_12_port, 
      position1_dp_cluster_4_add_178_aco_carry_13_port, 
      position1_dp_cluster_4_add_178_aco_carry_14_port, 
      position1_dp_cluster_4_add_178_aco_carry_15_port, 
      position1_dp_cluster_4_add_178_aco_carry_16_port, 
      position1_dp_cluster_4_add_178_aco_carry_17_port, 
      position1_dp_cluster_4_add_178_aco_carry_18_port, 
      position1_dp_cluster_4_add_178_aco_carry_19_port, 
      position1_dp_cluster_4_add_178_aco_carry_20_port, 
      position1_dp_cluster_4_add_178_aco_carry_21_port, 
      position1_dp_cluster_4_add_178_aco_carry_22_port, 
      position1_dp_cluster_4_add_178_aco_carry_23_port, 
      position1_dp_cluster_4_add_178_aco_carry_24_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_0_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_1_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_2_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_3_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_4_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_5_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_6_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_7_port, 
      position1_dp_cluster_5_mult_add_179_aco_PROD_not_8_port, 
      position1_dp_cluster_5_add_179_aco_carry_1_port, 
      position1_dp_cluster_5_add_179_aco_carry_2_port, 
      position1_dp_cluster_5_add_179_aco_carry_3_port, 
      position1_dp_cluster_5_add_179_aco_carry_4_port, 
      position1_dp_cluster_5_add_179_aco_carry_5_port, 
      position1_dp_cluster_5_add_179_aco_carry_6_port, 
      position1_dp_cluster_5_add_179_aco_carry_7_port, 
      position1_dp_cluster_5_add_179_aco_carry_8_port, 
      position1_dp_cluster_5_add_179_aco_carry_9_port, 
      position1_dp_cluster_5_add_179_aco_carry_10_port, 
      position1_dp_cluster_5_add_179_aco_carry_11_port, 
      position1_dp_cluster_5_add_179_aco_carry_12_port, 
      position1_dp_cluster_5_add_179_aco_carry_13_port, 
      position1_dp_cluster_5_add_179_aco_carry_14_port, 
      position1_dp_cluster_5_add_179_aco_carry_15_port, 
      position1_dp_cluster_5_add_179_aco_carry_16_port, 
      position1_dp_cluster_5_add_179_aco_carry_17_port, 
      position1_dp_cluster_5_add_179_aco_carry_18_port, 
      position1_dp_cluster_5_add_179_aco_carry_19_port, 
      position1_dp_cluster_5_add_179_aco_carry_20_port, 
      position1_dp_cluster_5_add_179_aco_carry_21_port, 
      position1_dp_cluster_5_add_179_aco_carry_22_port, 
      position1_dp_cluster_5_add_179_aco_carry_23_port, 
      position1_dp_cluster_5_add_179_aco_carry_24_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_2_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_3_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_4_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_5_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_6_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_7_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_8_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_9_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_10_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_11_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_12_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_13_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_14_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_15_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_16_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_17_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_18_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_19_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_20_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_21_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_22_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_23_port, 
      position1_dp_cluster_6_add_0_root_add_171_3_carry_24_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_2_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_3_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_4_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_5_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_6_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_7_port, 
      position1_dp_cluster_7_add_1_root_add_170_3_carry_8_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_2_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_3_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_4_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_5_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_6_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_7_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_8_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_9_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_10_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_11_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_12_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_13_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_14_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_15_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_16_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_17_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_18_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_19_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_20_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_21_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_22_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_23_port, 
      position1_dp_cluster_7_add_0_root_add_170_3_carry_24_port, 
      gensync1_add_39_carry_2_port, gensync1_add_39_carry_3_port, 
      gensync1_add_39_carry_4_port, gensync1_add_39_carry_5_port, 
      gensync1_add_39_carry_6_port, gensync1_add_39_carry_7_port, 
      gensync1_add_39_carry_8_port, gensync1_add_39_carry_9_port, 
      gensync1_add_45_carry_2_port, gensync1_add_45_carry_3_port, 
      gensync1_add_45_carry_4_port, gensync1_add_45_carry_5_port, 
      gensync1_add_45_carry_6_port, gensync1_add_45_carry_7_port, 
      gensync1_add_45_carry_8_port, gensync1_add_45_carry_9_port, 
      gensync1_sub_91_2_cf_carry_2_port, gensync1_sub_91_2_cf_carry_3_port, 
      gensync1_sub_91_2_cf_carry_4_port, gensync1_sub_91_2_cf_carry_5_port, 
      gensync1_sub_91_2_cf_carry_6_port, gensync1_sub_91_2_cf_carry_7_port, 
      gensync1_sub_91_2_cf_carry_8_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, 
      n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53
      , n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
      n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109
      , n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, cam_x_7_port,
      n493, cam_x_6_port, n495, cam_x_5_port, n497, cam_x_4_port, n499, 
      cam_x_3_port, n501, cam_x_2_port, n503, cam_x_1_port, n505, cam_x_0_port,
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, cam_y_0_port, IMG_top_port, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118 : std_logic;

begin
   r_out_proc <= ( r_out_proc_7_port, r_out_proc_6_port, r_out_proc_5_port, 
      r_out_proc_4_port, r_out_proc_3_port, r_out_proc_2_port, 
      r_out_proc_1_port, r_out_proc_0_port );
   g_out_proc <= ( g_out_proc_7_port, g_out_proc_6_port, g_out_proc_5_port, 
      g_out_proc_4_port, g_out_proc_3_port, g_out_proc_2_port, 
      g_out_proc_1_port, g_out_proc_0_port );
   b_out_proc <= ( b_out_proc_7_port, b_out_proc_6_port, b_out_proc_5_port, 
      b_out_proc_4_port, b_out_proc_3_port, b_out_proc_2_port, 
      b_out_proc_1_port, b_out_proc_0_port );
   X_barycentre_top <= ( X_barycentre_top_8_port, X_barycentre_top_7_port, 
      X_barycentre_top_6_port, X_barycentre_top_5_port, X_barycentre_top_4_port
      , X_barycentre_top_3_port, X_barycentre_top_2_port, 
      X_barycentre_top_1_port, X_barycentre_top_0_port );
   Y_barycentre_top <= ( Y_barycentre_top_8_port, Y_barycentre_top_7_port, 
      Y_barycentre_top_6_port, Y_barycentre_top_5_port, Y_barycentre_top_4_port
      , Y_barycentre_top_3_port, Y_barycentre_top_2_port, 
      Y_barycentre_top_1_port, Y_barycentre_top_0_port );
   cam_x <= ( cam_x_9_port, position1_dp_cluster_7_N314, cam_x_7_port, 
      cam_x_6_port, cam_x_5_port, cam_x_4_port, cam_x_3_port, cam_x_2_port, 
      cam_x_1_port, cam_x_0_port );
   cam_y <= ( position1_dp_cluster_6_N389, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, 
      position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, cam_y_0_port );
   IMG_top <= IMG_top_port;
   
   image_process1_U70 : OAI212 port map( A => n815, B => image_process1_n13, C 
                           => image_process1_n110, Q => image_process1_N14);
   image_process1_U68 : OAI212 port map( A => n815, B => image_process1_n25, C 
                           => image_process1_n110, Q => image_process1_N16);
   position1_U1019 : OAI212 port map( A => position1_N1519_port, B => n98, C =>
                           position1_n1578, Q => position1_N1573_port);
   position1_U1017 : OAI212 port map( A => position1_N1519_port, B => n92, C =>
                           position1_n1577, Q => position1_N1547_port);
   position1_U1015 : OAI212 port map( A => n520, B => n91, C => position1_n1576
                           , Q => position1_N1548_port);
   position1_U1013 : OAI212 port map( A => n522, B => n96, C => position1_n1575
                           , Q => position1_N1549_port);
   position1_U1011 : OAI212 port map( A => n522, B => n90, C => position1_n1574
                           , Q => position1_N1550_port);
   position1_U1009 : OAI212 port map( A => n522, B => n89, C => position1_n1573
                           , Q => position1_N1551_port);
   position1_U1007 : OAI212 port map( A => n522, B => n88, C => position1_n1572
                           , Q => position1_N1552_port);
   position1_U1005 : OAI212 port map( A => n522, B => n95, C => position1_n1571
                           , Q => position1_N1553_port);
   position1_U1003 : OAI212 port map( A => n522, B => n50, C => position1_n1570
                           , Q => position1_N1554_port);
   position1_U1001 : OAI212 port map( A => n522, B => n52, C => position1_n1569
                           , Q => position1_N1555_port);
   position1_U999 : OAI212 port map( A => n522, B => n70, C => position1_n1568,
                           Q => position1_N1556_port);
   position1_U997 : OAI212 port map( A => n522, B => n66, C => position1_n1567,
                           Q => position1_N1557_port);
   position1_U995 : OAI212 port map( A => n522, B => n82, C => position1_n1566,
                           Q => position1_N1558_port);
   position1_U993 : OAI212 port map( A => n522, B => n65, C => position1_n1565,
                           Q => position1_N1559_port);
   position1_U991 : OAI212 port map( A => n522, B => n81, C => position1_n1564,
                           Q => position1_N1560_port);
   position1_U989 : OAI212 port map( A => n522, B => n64, C => position1_n1563,
                           Q => position1_N1561_port);
   position1_U987 : OAI212 port map( A => n522, B => n80, C => position1_n1562,
                           Q => position1_N1562_port);
   position1_U985 : OAI212 port map( A => n522, B => n63, C => position1_n1561,
                           Q => position1_N1563_port);
   position1_U983 : OAI212 port map( A => n522, B => n79, C => position1_n1560,
                           Q => position1_N1564_port);
   position1_U981 : OAI212 port map( A => n521, B => n62, C => position1_n1559,
                           Q => position1_N1565_port);
   position1_U979 : OAI212 port map( A => n521, B => n78, C => position1_n1558,
                           Q => position1_N1566_port);
   position1_U977 : OAI212 port map( A => n520, B => n61, C => position1_n1557,
                           Q => position1_N1567_port);
   position1_U975 : OAI212 port map( A => position1_N1519_port, B => n77, C => 
                           position1_n1556, Q => position1_N1568_port);
   position1_U973 : OAI212 port map( A => position1_N1519_port, B => n60, C => 
                           position1_n1555, Q => position1_N1569_port);
   position1_U971 : OAI212 port map( A => position1_N1519_port, B => n100, C =>
                           position1_n1554, Q => position1_N1570_port);
   position1_U945 : OAI222 port map( A => n530, B => position1_n1553, C => n528
                           , D => position1_n1553, Q => position1_N1677);
   position1_U944 : OAI222 port map( A => n531, B => position1_n1552, C => n528
                           , D => position1_n1552, Q => position1_N1651);
   position1_U943 : OAI222 port map( A => n531, B => position1_n1551, C => n528
                           , D => position1_n1551, Q => position1_N1652);
   position1_U942 : OAI222 port map( A => n531, B => position1_n1550, C => n528
                           , D => position1_n1550, Q => position1_N1653);
   position1_U941 : OAI222 port map( A => n531, B => position1_n1549, C => n528
                           , D => position1_n1549, Q => position1_N1654);
   position1_U940 : OAI222 port map( A => n531, B => position1_n1548, C => n528
                           , D => position1_n1548, Q => position1_N1655);
   position1_U939 : OAI222 port map( A => n531, B => n105, C => n528, D => 
                           position1_n1547, Q => position1_N1656);
   position1_U938 : OAI222 port map( A => n531, B => n1299, C => n528, D => 
                           position1_n1546, Q => position1_N1657);
   position1_U937 : OAI222 port map( A => n531, B => n1296, C => n528, D => 
                           position1_n1545, Q => position1_N1658);
   position1_U936 : OAI222 port map( A => n531, B => n1294, C => n528, D => 
                           position1_n1544, Q => position1_N1659);
   position1_U935 : OAI222 port map( A => n531, B => n1291, C => n528, D => 
                           position1_n1543, Q => position1_N1660);
   position1_U934 : OAI222 port map( A => n532, B => n1289, C => n528, D => 
                           position1_n1542, Q => position1_N1661);
   position1_U933 : OAI222 port map( A => n532, B => n1287, C => n528, D => 
                           position1_n1541, Q => position1_N1662);
   position1_U932 : OAI222 port map( A => n532, B => n1285, C => n529, D => 
                           position1_n1540, Q => position1_N1663);
   position1_U931 : OAI222 port map( A => n532, B => n1283, C => n529, D => 
                           position1_n1539, Q => position1_N1664);
   position1_U930 : OAI222 port map( A => n530, B => n1281, C => n529, D => 
                           position1_n1538, Q => position1_N1665);
   position1_U929 : OAI222 port map( A => n532, B => n1279, C => n529, D => 
                           position1_n1537, Q => position1_N1666);
   position1_U928 : OAI222 port map( A => n530, B => n1277, C => n529, D => 
                           position1_n1536, Q => position1_N1667);
   position1_U927 : OAI222 port map( A => n532, B => n1275, C => n529, D => 
                           position1_n1535, Q => position1_N1668);
   position1_U926 : OAI222 port map( A => n532, B => n1273, C => n529, D => 
                           position1_n1534, Q => position1_N1669);
   position1_U925 : OAI222 port map( A => n532, B => n1271, C => n529, D => 
                           position1_n1533, Q => position1_N1670);
   position1_U924 : OAI222 port map( A => n530, B => n1250, C => n529, D => 
                           position1_n1532, Q => position1_N1671);
   position1_U923 : OAI222 port map( A => n530, B => n1248, C => n529, D => 
                           position1_n1531, Q => position1_N1672);
   position1_U922 : OAI222 port map( A => n530, B => n1247, C => n529, D => 
                           position1_n1530, Q => position1_N1673);
   position1_U921 : OAI222 port map( A => n530, B => n107, C => n529, D => 
                           position1_n1529, Q => position1_N1674);
   position1_U799 : OAI212 port map( A => position1_state_1_port, B => 
                           position1_state_0_port, C => n488, Q => 
                           position1_N2353);
   position1_U783 : OAI212 port map( A => position1_n1395, B => position1_n1396
                           , C => n853, Q => position1_n1390);
   position1_U773 : OAI222 port map( A => n1360, B => n654, C => 
                           position1_n1141, D => position1_n1064, Q => 
                           position1_N193);
   position1_U764 : OAI212 port map( A => position1_N1936, B => n97, C => 
                           position1_n1382, Q => position1_N1990);
   position1_U762 : OAI212 port map( A => position1_N1936, B => n87, C => 
                           position1_n1381, Q => position1_N1964);
   position1_U760 : OAI212 port map( A => n554, B => n86, C => position1_n1380,
                           Q => position1_N1965);
   position1_U758 : OAI212 port map( A => n556, B => n94, C => position1_n1379,
                           Q => position1_N1966);
   position1_U756 : OAI212 port map( A => n556, B => n85, C => position1_n1378,
                           Q => position1_N1967);
   position1_U754 : OAI212 port map( A => n556, B => n84, C => position1_n1377,
                           Q => position1_N1968);
   position1_U752 : OAI212 port map( A => n556, B => n83, C => position1_n1376,
                           Q => position1_N1969);
   position1_U750 : OAI212 port map( A => n556, B => n93, C => position1_n1375,
                           Q => position1_N1970);
   position1_U748 : OAI212 port map( A => n556, B => n49, C => position1_n1374,
                           Q => position1_N1971);
   position1_U746 : OAI212 port map( A => n556, B => n51, C => position1_n1373,
                           Q => position1_N1972);
   position1_U744 : OAI212 port map( A => n556, B => n69, C => position1_n1372,
                           Q => position1_N1973);
   position1_U742 : OAI212 port map( A => n556, B => n59, C => position1_n1371,
                           Q => position1_N1974);
   position1_U740 : OAI212 port map( A => n556, B => n76, C => position1_n1370,
                           Q => position1_N1975);
   position1_U738 : OAI212 port map( A => n556, B => n58, C => position1_n1369,
                           Q => position1_N1976);
   position1_U736 : OAI212 port map( A => n556, B => n75, C => position1_n1368,
                           Q => position1_N1977);
   position1_U734 : OAI212 port map( A => n556, B => n57, C => position1_n1367,
                           Q => position1_N1978);
   position1_U732 : OAI212 port map( A => n556, B => n74, C => position1_n1366,
                           Q => position1_N1979);
   position1_U730 : OAI212 port map( A => n556, B => n56, C => position1_n1365,
                           Q => position1_N1980);
   position1_U728 : OAI212 port map( A => n556, B => n73, C => position1_n1364,
                           Q => position1_N1981);
   position1_U726 : OAI212 port map( A => n555, B => n55, C => position1_n1363,
                           Q => position1_N1982);
   position1_U724 : OAI212 port map( A => n555, B => n72, C => position1_n1362,
                           Q => position1_N1983);
   position1_U722 : OAI212 port map( A => n554, B => n54, C => position1_n1361,
                           Q => position1_N1984);
   position1_U720 : OAI212 port map( A => position1_N1936, B => n71, C => 
                           position1_n1360, Q => position1_N1985);
   position1_U718 : OAI212 port map( A => position1_N1936, B => n53, C => 
                           position1_n1359, Q => position1_N1986);
   position1_U716 : OAI212 port map( A => position1_N1936, B => n99, C => 
                           position1_n1358, Q => position1_N1987);
   position1_U690 : OAI222 port map( A => n564, B => position1_n1357, C => n562
                           , D => position1_n1357, Q => position1_N2094);
   position1_U689 : OAI222 port map( A => n565, B => position1_n1356, C => n562
                           , D => position1_n1356, Q => position1_N2068);
   position1_U688 : OAI222 port map( A => n565, B => position1_n1355, C => n562
                           , D => position1_n1355, Q => position1_N2069);
   position1_U687 : OAI222 port map( A => n565, B => position1_n1354, C => n562
                           , D => position1_n1354, Q => position1_N2070);
   position1_U686 : OAI222 port map( A => n565, B => position1_n1353, C => n562
                           , D => position1_n1353, Q => position1_N2071);
   position1_U685 : OAI222 port map( A => n565, B => position1_n1352, C => n562
                           , D => position1_n1352, Q => position1_N2072);
   position1_U684 : OAI222 port map( A => n565, B => n106, C => n562, D => 
                           position1_n1351, Q => position1_N2073);
   position1_U683 : OAI222 port map( A => n565, B => n1080, C => n562, D => 
                           position1_n1350, Q => position1_N2074);
   position1_U682 : OAI222 port map( A => n565, B => n1077, C => n562, D => 
                           position1_n1349, Q => position1_N2075);
   position1_U681 : OAI222 port map( A => n565, B => n1075, C => n562, D => 
                           position1_n1348, Q => position1_N2076);
   position1_U680 : OAI222 port map( A => n565, B => n1072, C => n562, D => 
                           position1_n1347, Q => position1_N2077);
   position1_U679 : OAI222 port map( A => n566, B => n1070, C => n562, D => 
                           position1_n1346, Q => position1_N2078);
   position1_U678 : OAI222 port map( A => n566, B => n1068, C => n562, D => 
                           position1_n1345, Q => position1_N2079);
   position1_U677 : OAI222 port map( A => n566, B => n1066, C => n563, D => 
                           position1_n1344, Q => position1_N2080);
   position1_U676 : OAI222 port map( A => n566, B => n1064, C => n563, D => 
                           position1_n1343, Q => position1_N2081);
   position1_U675 : OAI222 port map( A => n564, B => n1062, C => n563, D => 
                           position1_n1342, Q => position1_N2082);
   position1_U674 : OAI222 port map( A => n566, B => n1060, C => n563, D => 
                           position1_n1341, Q => position1_N2083);
   position1_U673 : OAI222 port map( A => n564, B => n1058, C => n563, D => 
                           position1_n1340, Q => position1_N2084);
   position1_U672 : OAI222 port map( A => n566, B => n1056, C => n563, D => 
                           position1_n1339, Q => position1_N2085);
   position1_U671 : OAI222 port map( A => n566, B => n1054, C => n563, D => 
                           position1_n1338, Q => position1_N2086);
   position1_U670 : OAI222 port map( A => n566, B => n1052, C => n563, D => 
                           position1_n1337, Q => position1_N2087);
   position1_U669 : OAI222 port map( A => n564, B => n1031, C => n563, D => 
                           position1_n1336, Q => position1_N2088);
   position1_U668 : OAI222 port map( A => n564, B => n1029, C => n563, D => 
                           position1_n1335, Q => position1_N2089);
   position1_U667 : OAI222 port map( A => n564, B => n1028, C => n563, D => 
                           position1_n1334, Q => position1_N2090);
   position1_U666 : OAI222 port map( A => n564, B => n108, C => n563, D => 
                           position1_n1333, Q => position1_N2091);
   position1_U487 : OAI212 port map( A => n656, B => position1_n362, C => n714,
                           Q => position1_N89);
   position1_U485 : OAI212 port map( A => n656, B => position1_n360, C => n714,
                           Q => position1_N91);
   position1_U483 : OAI212 port map( A => n655, B => position1_n358, C => n714,
                           Q => position1_N93);
   position1_U482 : OAI212 port map( A => n654, B => position1_n357, C => n714,
                           Q => position1_N94);
   position1_U481 : OAI212 port map( A => n654, B => position1_n356, C => n714,
                           Q => position1_N95);
   position1_U447 : OAI222 port map( A => position1_n1063, B => position1_n1151
                           , C => position1_n1141, D => position1_n1145, Q => 
                           position1_n1072);
   position1_U445 : OAI222 port map( A => position1_n1149, B => position1_n1062
                           , C => position1_n1146, D => position1_n1141, Q => 
                           position1_n1060);
   position1_U438 : OAI222 port map( A => position1_n1062, B => position1_n1065
                           , C => position1_n1141, D => position1_n1058, Q => 
                           position1_n1071);
   position1_r406_U1_1 : ADD32 port map( A => position1_x_sum_1_port, B => 
                           cam_x_1_port, CI => position1_r406_carry_1_port, CO 
                           => position1_r406_carry_2_port, S => position1_N281)
                           ;
   position1_r406_U1_2 : ADD32 port map( A => position1_x_sum_2_port, B => 
                           cam_x_2_port, CI => position1_r406_carry_2_port, CO 
                           => position1_r406_carry_3_port, S => position1_N282)
                           ;
   position1_r406_U1_3 : ADD32 port map( A => position1_x_sum_3_port, B => 
                           cam_x_3_port, CI => position1_r406_carry_3_port, CO 
                           => position1_r406_carry_4_port, S => 
                           position1_N283_port);
   position1_r406_U1_4 : ADD32 port map( A => position1_x_sum_4_port, B => 
                           cam_x_4_port, CI => position1_r406_carry_4_port, CO 
                           => position1_r406_carry_5_port, S => position1_N284)
                           ;
   position1_r406_U1_5 : ADD32 port map( A => position1_x_sum_5_port, B => 
                           cam_x_5_port, CI => position1_r406_carry_5_port, CO 
                           => position1_r406_carry_6_port, S => position1_N285)
                           ;
   position1_r406_U1_6 : ADD32 port map( A => position1_x_sum_6_port, B => 
                           cam_x_6_port, CI => position1_r406_carry_6_port, CO 
                           => position1_r406_carry_7_port, S => position1_N286)
                           ;
   position1_r406_U1_7 : ADD32 port map( A => position1_x_sum_7_port, B => 
                           cam_x_7_port, CI => position1_r406_carry_7_port, CO 
                           => position1_r406_carry_8_port, S => position1_N287)
                           ;
   position1_r406_U1_8 : ADD32 port map( A => position1_x_sum_8_port, B => 
                           position1_dp_cluster_7_N314, CI => 
                           position1_r406_carry_8_port, CO => 
                           position1_r406_carry_9_port, S => position1_N288);
   position1_r409_U1_1 : ADD32 port map( A => position1_y_sum_1_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, 
                           CI => position1_r409_carry_1_port, CO => 
                           position1_r409_carry_2_port, S => 
                           position1_N356_port);
   position1_r409_U1_2 : ADD32 port map( A => position1_y_sum_2_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, 
                           CI => position1_r409_carry_2_port, CO => 
                           position1_r409_carry_3_port, S => 
                           position1_N357_port);
   position1_r409_U1_3 : ADD32 port map( A => position1_y_sum_3_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, 
                           CI => position1_r409_carry_3_port, CO => 
                           position1_r409_carry_4_port, S => 
                           position1_N358_port);
   position1_r409_U1_4 : ADD32 port map( A => position1_y_sum_4_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, 
                           CI => position1_r409_carry_4_port, CO => 
                           position1_r409_carry_5_port, S => position1_N359);
   position1_r409_U1_5 : ADD32 port map( A => position1_y_sum_5_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, 
                           CI => position1_r409_carry_5_port, CO => 
                           position1_r409_carry_6_port, S => 
                           position1_N360_port);
   position1_r409_U1_6 : ADD32 port map( A => position1_y_sum_6_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, 
                           CI => position1_r409_carry_6_port, CO => 
                           position1_r409_carry_7_port, S => position1_N361);
   position1_r409_U1_7 : ADD32 port map( A => position1_y_sum_7_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, 
                           CI => position1_r409_carry_7_port, CO => 
                           position1_r409_carry_8_port, S => 
                           position1_N362_port);
   position1_r409_U1_8 : ADD32 port map( A => position1_y_sum_8_port, B => 
                           position1_dp_cluster_6_N389, CI => 
                           position1_r409_carry_8_port, CO => 
                           position1_r409_carry_9_port, S => 
                           position1_N363_port);
   position1_r412_U1_1 : ADD32 port map( A => n503, B => position1_N281, CI => 
                           position1_r412_carry_1_port, CO => 
                           position1_r412_carry_2_port, S => position1_N486);
   position1_r412_U1_2 : ADD32 port map( A => n501, B => position1_N282, CI => 
                           position1_r412_carry_2_port, CO => 
                           position1_r412_carry_3_port, S => position1_N487);
   position1_r412_U1_3 : ADD32 port map( A => n499, B => position1_N283_port, 
                           CI => position1_r412_carry_3_port, CO => 
                           position1_r412_carry_4_port, S => position1_N488);
   position1_r412_U1_4 : ADD32 port map( A => n497, B => position1_N284, CI => 
                           position1_r412_carry_4_port, CO => 
                           position1_r412_carry_5_port, S => position1_N489);
   position1_r412_U1_5 : ADD32 port map( A => n495, B => position1_N285, CI => 
                           position1_r412_carry_5_port, CO => 
                           position1_r412_carry_6_port, S => position1_N490);
   position1_r412_U1_6 : ADD32 port map( A => n493, B => position1_N286, CI => 
                           position1_r412_carry_6_port, CO => 
                           position1_r412_carry_7_port, S => position1_N491);
   position1_r412_U1_7 : ADD32 port map( A => n491, B => position1_N287, CI => 
                           position1_r412_carry_7_port, CO => 
                           position1_r412_carry_8_port, S => position1_N492);
   position1_r412_U1_8 : ADD32 port map( A => position1_dp_cluster_7_N314, B =>
                           position1_N288, CI => position1_r412_carry_8_port, 
                           CO => position1_r412_carry_9_port, S => 
                           position1_N493);
   position1_r413_U1_1 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, B 
                           => position1_N356_port, CI => 
                           position1_r413_carry_1_port, CO => 
                           position1_r413_carry_2_port, S => position1_N536);
   position1_r413_U1_2 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, B 
                           => position1_N357_port, CI => 
                           position1_r413_carry_2_port, CO => 
                           position1_r413_carry_3_port, S => position1_N537);
   position1_r413_U1_3 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => position1_N358_port, CI => 
                           position1_r413_carry_3_port, CO => 
                           position1_r413_carry_4_port, S => position1_N538);
   position1_r413_U1_4 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, B 
                           => position1_N359, CI => position1_r413_carry_4_port
                           , CO => position1_r413_carry_5_port, S => 
                           position1_N539);
   position1_r413_U1_5 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, B 
                           => position1_N360_port, CI => 
                           position1_r413_carry_5_port, CO => 
                           position1_r413_carry_6_port, S => position1_N540);
   position1_r413_U1_6 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, B 
                           => position1_N361, CI => position1_r413_carry_6_port
                           , CO => position1_r413_carry_7_port, S => 
                           position1_N541);
   position1_r413_U1_7 : ADD32 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, B 
                           => position1_N362_port, CI => 
                           position1_r413_carry_7_port, CO => 
                           position1_r413_carry_8_port, S => position1_N542);
   position1_r413_U1_8 : ADD32 port map( A => position1_dp_cluster_6_N389, B =>
                           position1_N363_port, CI => 
                           position1_r413_carry_8_port, CO => 
                           position1_r413_carry_9_port, S => position1_N543);
   position1_r416_U1_1_1 : ADD22 port map( A => n633, B => n516, CO => 
                           position1_r416_carry_2_port, S => position1_N590);
   position1_r416_U1_1_2 : ADD22 port map( A => n629, B => 
                           position1_r416_carry_2_port, CO => 
                           position1_r416_carry_3_port, S => position1_N591);
   position1_r416_U1_1_3 : ADD22 port map( A => n625, B => 
                           position1_r416_carry_3_port, CO => 
                           position1_r416_carry_4_port, S => position1_N592);
   position1_r416_U1_1_4 : ADD22 port map( A => n469, B => 
                           position1_r416_carry_4_port, CO => 
                           position1_r416_carry_5_port, S => position1_N593);
   position1_r416_U1_1_5 : ADD22 port map( A => n622, B => 
                           position1_r416_carry_5_port, CO => 
                           position1_r416_carry_6_port, S => position1_N594);
   position1_r416_U1_1_6 : ADD22 port map( A => n470, B => 
                           position1_r416_carry_6_port, CO => 
                           position1_r416_carry_7_port, S => position1_N595);
   position1_r416_U1_1_7 : ADD22 port map( A => n617, B => 
                           position1_r416_carry_7_port, CO => 
                           position1_r416_carry_8_port, S => position1_N596);
   position1_r416_U1_1_8 : ADD22 port map( A => n472, B => 
                           position1_r416_carry_8_port, CO => 
                           position1_r416_carry_9_port, S => position1_N597);
   position1_r416_U1_1_9 : ADD22 port map( A => n610, B => 
                           position1_r416_carry_9_port, CO => 
                           position1_r416_carry_10_port, S => position1_N598);
   position1_r416_U1_1_10 : ADD22 port map( A => n474, B => 
                           position1_r416_carry_10_port, CO => 
                           position1_r416_carry_11_port, S => position1_N599);
   position1_r416_U1_1_11 : ADD22 port map( A => n607, B => 
                           position1_r416_carry_11_port, CO => 
                           position1_r416_carry_12_port, S => position1_N600);
   position1_r416_U1_1_12 : ADD22 port map( A => n475, B => 
                           position1_r416_carry_12_port, CO => 
                           position1_r416_carry_13_port, S => position1_N601);
   position1_r416_U1_1_13 : ADD22 port map( A => n603, B => 
                           position1_r416_carry_13_port, CO => 
                           position1_r416_carry_14_port, S => position1_N602);
   position1_r416_U1_1_14 : ADD22 port map( A => n476, B => 
                           position1_r416_carry_14_port, CO => 
                           position1_r416_carry_15_port, S => position1_N603);
   position1_r416_U1_1_15 : ADD22 port map( A => n599, B => 
                           position1_r416_carry_15_port, CO => 
                           position1_r416_carry_16_port, S => position1_N604);
   position1_r416_U1_1_16 : ADD22 port map( A => n596, B => 
                           position1_r416_carry_16_port, CO => 
                           position1_r416_carry_17_port, S => position1_N605);
   position1_add_161_U1_1_1 : ADD22 port map( A => position1_count_img_1_port, 
                           B => position1_count_img_0_port, CO => 
                           position1_add_161_carry_2_port, S => position1_N206)
                           ;
   position1_add_161_U1_1_2 : ADD22 port map( A => position1_count_img_2_port, 
                           B => position1_add_161_carry_2_port, CO => 
                           position1_add_161_carry_3_port, S => position1_N207)
                           ;
   position1_add_161_U1_1_3 : ADD22 port map( A => position1_count_img_3_port, 
                           B => position1_add_161_carry_3_port, CO => 
                           position1_add_161_carry_4_port, S => position1_N208)
                           ;
   position1_add_161_U1_1_4 : ADD22 port map( A => position1_count_img_4_port, 
                           B => position1_add_161_carry_4_port, CO => 
                           position1_add_161_carry_5_port, S => position1_N209)
                           ;
   position1_add_161_U1_1_5 : ADD22 port map( A => position1_count_img_5_port, 
                           B => position1_add_161_carry_5_port, CO => 
                           position1_add_161_carry_6_port, S => position1_N210)
                           ;
   position1_add_161_U1_1_6 : ADD22 port map( A => position1_count_img_6_port, 
                           B => position1_add_161_carry_6_port, CO => 
                           position1_add_161_carry_7_port, S => position1_N211)
                           ;
   position1_add_161_U1_1_7 : ADD22 port map( A => position1_count_img_7_port, 
                           B => position1_add_161_carry_7_port, CO => 
                           position1_add_161_carry_8_port, S => position1_N212)
                           ;
   position1_add_161_U1_1_8 : ADD22 port map( A => position1_count_img_8_port, 
                           B => position1_add_161_carry_8_port, CO => 
                           position1_add_161_carry_9_port, S => position1_N213)
                           ;
   position1_add_161_U1_1_9 : ADD22 port map( A => position1_count_img_9_port, 
                           B => position1_add_161_carry_9_port, CO => 
                           position1_add_161_carry_10_port, S => position1_N214
                           );
   position1_add_161_U1_1_10 : ADD22 port map( A => position1_count_img_10_port
                           , B => position1_add_161_carry_10_port, CO => 
                           position1_add_161_carry_11_port, S => position1_N215
                           );
   position1_add_161_U1_1_11 : ADD22 port map( A => position1_count_img_11_port
                           , B => position1_add_161_carry_11_port, CO => 
                           position1_add_161_carry_12_port, S => position1_N216
                           );
   position1_add_161_U1_1_12 : ADD22 port map( A => position1_count_img_12_port
                           , B => position1_add_161_carry_12_port, CO => 
                           position1_add_161_carry_13_port, S => position1_N217
                           );
   position1_add_161_U1_1_13 : ADD22 port map( A => position1_count_img_13_port
                           , B => position1_add_161_carry_13_port, CO => 
                           position1_add_161_carry_14_port, S => position1_N218
                           );
   position1_add_161_U1_1_14 : ADD22 port map( A => position1_count_img_14_port
                           , B => position1_add_161_carry_14_port, CO => 
                           position1_add_161_carry_15_port, S => position1_N219
                           );
   position1_add_161_U1_1_15 : ADD22 port map( A => position1_count_img_15_port
                           , B => position1_add_161_carry_15_port, CO => 
                           position1_add_161_carry_16_port, S => position1_N220
                           );
   position1_add_161_U1_1_16 : ADD22 port map( A => position1_count_img_16_port
                           , B => position1_add_161_carry_16_port, CO => 
                           position1_add_161_carry_17_port, S => position1_N221
                           );
   position1_add_161_U1_1_17 : ADD22 port map( A => position1_count_img_17_port
                           , B => position1_add_161_carry_17_port, CO => 
                           position1_add_161_carry_18_port, S => position1_N222
                           );
   position1_add_161_U1_1_18 : ADD22 port map( A => position1_count_img_18_port
                           , B => position1_add_161_carry_18_port, CO => 
                           position1_add_161_carry_19_port, S => position1_N223
                           );
   position1_sub_216_U2_9 : ADD32 port map( A => position1_x_sum_9_port, B => 
                           n630, CI => position1_sub_216_carry_9_port, CO => 
                           position1_sub_216_carry_10_port, S => 
                           position1_N1530_port);
   position1_sub_216_U2_10 : ADD32 port map( A => position1_x_sum_10_port, B =>
                           n67, CI => position1_sub_216_carry_10_port, CO => 
                           position1_sub_216_carry_11_port, S => 
                           position1_N1531_port);
   position1_sub_216_U2_11 : ADD32 port map( A => position1_x_sum_11_port, B =>
                           n274, CI => position1_sub_216_carry_11_port, CO => 
                           position1_sub_216_carry_12_port, S => 
                           position1_N1532_port);
   position1_sub_216_U2_12 : ADD32 port map( A => position1_x_sum_12_port, B =>
                           n42, CI => position1_sub_216_carry_12_port, CO => 
                           position1_sub_216_carry_13_port, S => 
                           position1_N1533_port);
   position1_sub_216_U2_13 : ADD32 port map( A => position1_x_sum_13_port, B =>
                           n278, CI => position1_sub_216_carry_13_port, CO => 
                           position1_sub_216_carry_14_port, S => 
                           position1_N1534_port);
   position1_sub_216_U2_14 : ADD32 port map( A => position1_x_sum_14_port, B =>
                           n280, CI => position1_sub_216_carry_14_port, CO => 
                           position1_sub_216_carry_15_port, S => 
                           position1_N1535_port);
   position1_sub_216_U2_15 : ADD32 port map( A => position1_x_sum_15_port, B =>
                           n282, CI => position1_sub_216_carry_15_port, CO => 
                           position1_sub_216_carry_16_port, S => 
                           position1_N1536_port);
   position1_sub_216_U2_16 : ADD32 port map( A => position1_x_sum_16_port, B =>
                           n41, CI => position1_sub_216_carry_16_port, CO => 
                           position1_sub_216_carry_17_port, S => 
                           position1_N1537_port);
   position1_sub_216_U2_17 : ADD32 port map( A => position1_x_sum_17_port, B =>
                           n286, CI => position1_sub_216_carry_17_port, CO => 
                           position1_sub_216_carry_18_port, S => 
                           position1_N1538_port);
   position1_sub_216_U2_18 : ADD32 port map( A => position1_x_sum_18_port, B =>
                           n47, CI => position1_sub_216_carry_18_port, CO => 
                           position1_sub_216_carry_19_port, S => 
                           position1_N1539_port);
   position1_sub_216_U2_19 : ADD32 port map( A => position1_x_sum_19_port, B =>
                           n290, CI => position1_sub_216_carry_19_port, CO => 
                           position1_sub_216_carry_20_port, S => 
                           position1_N1540_port);
   position1_sub_216_U2_20 : ADD32 port map( A => position1_x_sum_20_port, B =>
                           n44, CI => position1_sub_216_carry_20_port, CO => 
                           position1_sub_216_carry_21_port, S => 
                           position1_N1541_port);
   position1_sub_216_U2_21 : ADD32 port map( A => position1_x_sum_21_port, B =>
                           n294, CI => position1_sub_216_carry_21_port, CO => 
                           position1_sub_216_carry_22_port, S => 
                           position1_N1542_port);
   position1_sub_216_U2_22 : ADD32 port map( A => position1_x_sum_22_port, B =>
                           n43, CI => position1_sub_216_carry_22_port, CO => 
                           position1_sub_216_carry_23_port, S => 
                           position1_N1543_port);
   position1_sub_216_U2_23 : ADD32 port map( A => position1_x_sum_23_port, B =>
                           n298, CI => position1_sub_216_carry_23_port, CO => 
                           position1_sub_216_carry_24_port, S => 
                           position1_N1544_port);
   position1_sub_216_I2_U2_8 : ADD32 port map( A => position1_N1554_port, B => 
                           n37, CI => position1_sub_216_I2_carry_8_port, CO => 
                           position1_sub_216_I2_carry_9_port, S => 
                           position1_N1581_port);
   position1_sub_216_I2_U2_9 : ADD32 port map( A => position1_N1555_port, B => 
                           n272, CI => position1_sub_216_I2_carry_9_port, CO =>
                           position1_sub_216_I2_carry_10_port, S => 
                           position1_N1582_port);
   position1_sub_216_I2_U2_10 : ADD32 port map( A => position1_N1556_port, B =>
                           n274, CI => position1_sub_216_I2_carry_10_port, CO 
                           => position1_sub_216_I2_carry_11_port, S => 
                           position1_N1583_port);
   position1_sub_216_I2_U2_11 : ADD32 port map( A => position1_N1557_port, B =>
                           n276, CI => position1_sub_216_I2_carry_11_port, CO 
                           => position1_sub_216_I2_carry_12_port, S => 
                           position1_N1584_port);
   position1_sub_216_I2_U2_12 : ADD32 port map( A => position1_N1558_port, B =>
                           n278, CI => position1_sub_216_I2_carry_12_port, CO 
                           => position1_sub_216_I2_carry_13_port, S => 
                           position1_N1585_port);
   position1_sub_216_I2_U2_13 : ADD32 port map( A => position1_N1559_port, B =>
                           n280, CI => position1_sub_216_I2_carry_13_port, CO 
                           => position1_sub_216_I2_carry_14_port, S => 
                           position1_N1586_port);
   position1_sub_216_I2_U2_14 : ADD32 port map( A => position1_N1560_port, B =>
                           n282, CI => position1_sub_216_I2_carry_14_port, CO 
                           => position1_sub_216_I2_carry_15_port, S => 
                           position1_N1587_port);
   position1_sub_216_I2_U2_15 : ADD32 port map( A => position1_N1561_port, B =>
                           n256, CI => position1_sub_216_I2_carry_15_port, CO 
                           => position1_sub_216_I2_carry_16_port, S => 
                           position1_N1588_port);
   position1_sub_216_I2_U2_16 : ADD32 port map( A => position1_N1562_port, B =>
                           n36, CI => position1_sub_216_I2_carry_16_port, CO =>
                           position1_sub_216_I2_carry_17_port, S => 
                           position1_N1589_port);
   position1_sub_216_I2_U2_17 : ADD32 port map( A => position1_N1563_port, B =>
                           n288, CI => position1_sub_216_I2_carry_17_port, CO 
                           => position1_sub_216_I2_carry_18_port, S => 
                           position1_N1590_port);
   position1_sub_216_I2_U2_18 : ADD32 port map( A => position1_N1564_port, B =>
                           n290, CI => position1_sub_216_I2_carry_18_port, CO 
                           => position1_sub_216_I2_carry_19_port, S => 
                           position1_N1591_port);
   position1_sub_216_I2_U2_19 : ADD32 port map( A => position1_N1565_port, B =>
                           n263, CI => position1_sub_216_I2_carry_19_port, CO 
                           => position1_sub_216_I2_carry_20_port, S => 
                           position1_N1592_port);
   position1_sub_216_I2_U2_20 : ADD32 port map( A => position1_N1566_port, B =>
                           n294, CI => position1_sub_216_I2_carry_20_port, CO 
                           => position1_sub_216_I2_carry_21_port, S => 
                           position1_N1593_port);
   position1_sub_216_I2_U2_21 : ADD32 port map( A => position1_N1567_port, B =>
                           n296, CI => position1_sub_216_I2_carry_21_port, CO 
                           => position1_sub_216_I2_carry_22_port, S => 
                           position1_N1594_port);
   position1_sub_216_I2_U2_22 : ADD32 port map( A => position1_N1568_port, B =>
                           n269, CI => position1_sub_216_I2_carry_22_port, CO 
                           => position1_sub_216_I2_carry_23_port, S => 
                           position1_N1595_port);
   position1_sub_216_I2_U2_23 : ADD32 port map( A => position1_N1569_port, B =>
                           n300, CI => position1_sub_216_I2_carry_23_port, CO 
                           => position1_sub_216_I2_carry_24_port, S => 
                           position1_N1596_port);
   position1_sub_216_I3_U2_7 : ADD32 port map( A => n1300, B => n37, CI => 
                           position1_sub_216_I3_carry_7_port, CO => 
                           position1_sub_216_I3_carry_8_port, S => 
                           position1_N1632_port);
   position1_sub_216_I3_U2_8 : ADD32 port map( A => n1298, B => n245, CI => 
                           position1_sub_216_I3_carry_8_port, CO => 
                           position1_sub_216_I3_carry_9_port, S => 
                           position1_N1633_port);
   position1_sub_216_I3_U2_9 : ADD32 port map( A => n1295, B => n246, CI => 
                           position1_sub_216_I3_carry_9_port, CO => 
                           position1_sub_216_I3_carry_10_port, S => 
                           position1_N1634_port);
   position1_sub_216_I3_U2_10 : ADD32 port map( A => n1293, B => n248, CI => 
                           position1_sub_216_I3_carry_10_port, CO => 
                           position1_sub_216_I3_carry_11_port, S => 
                           position1_N1635_port);
   position1_sub_216_I3_U2_11 : ADD32 port map( A => n1290, B => n48, CI => 
                           position1_sub_216_I3_carry_11_port, CO => 
                           position1_sub_216_I3_carry_12_port, S => 
                           position1_N1636);
   position1_sub_216_I3_U2_12 : ADD32 port map( A => n1288, B => n252, CI => 
                           position1_sub_216_I3_carry_12_port, CO => 
                           position1_sub_216_I3_carry_13_port, S => 
                           position1_N1637);
   position1_sub_216_I3_U2_13 : ADD32 port map( A => n1286, B => n254, CI => 
                           position1_sub_216_I3_carry_13_port, CO => 
                           position1_sub_216_I3_carry_14_port, S => 
                           position1_N1638);
   position1_sub_216_I3_U2_14 : ADD32 port map( A => n1284, B => n284, CI => 
                           position1_sub_216_I3_carry_14_port, CO => 
                           position1_sub_216_I3_carry_15_port, S => 
                           position1_N1639);
   position1_sub_216_I3_U2_15 : ADD32 port map( A => n1282, B => n286, CI => 
                           position1_sub_216_I3_carry_15_port, CO => 
                           position1_sub_216_I3_carry_16_port, S => 
                           position1_N1640);
   position1_sub_216_I3_U2_16 : ADD32 port map( A => n1280, B => n259, CI => 
                           position1_sub_216_I3_carry_16_port, CO => 
                           position1_sub_216_I3_carry_17_port, S => 
                           position1_N1641);
   position1_sub_216_I3_U2_17 : ADD32 port map( A => n1278, B => n261, CI => 
                           position1_sub_216_I3_carry_17_port, CO => 
                           position1_sub_216_I3_carry_18_port, S => 
                           position1_N1642);
   position1_sub_216_I3_U2_18 : ADD32 port map( A => n1276, B => n292, CI => 
                           position1_sub_216_I3_carry_18_port, CO => 
                           position1_sub_216_I3_carry_19_port, S => 
                           position1_N1643);
   position1_sub_216_I3_U2_19 : ADD32 port map( A => n1274, B => n265, CI => 
                           position1_sub_216_I3_carry_19_port, CO => 
                           position1_sub_216_I3_carry_20_port, S => 
                           position1_N1644);
   position1_sub_216_I3_U2_20 : ADD32 port map( A => n1272, B => n267, CI => 
                           position1_sub_216_I3_carry_20_port, CO => 
                           position1_sub_216_I3_carry_21_port, S => 
                           position1_N1645);
   position1_sub_216_I3_U2_21 : ADD32 port map( A => n1270, B => n68, CI => 
                           position1_sub_216_I3_carry_21_port, CO => 
                           position1_sub_216_I3_carry_22_port, S => 
                           position1_N1646);
   position1_sub_216_I3_U2_22 : ADD32 port map( A => n1269, B => n45, CI => 
                           position1_sub_216_I3_carry_22_port, CO => 
                           position1_sub_216_I3_carry_23_port, S => 
                           position1_N1647);
   position1_sub_216_I3_U2_23 : ADD32 port map( A => n1268, B => n589, CI => 
                           position1_sub_216_I3_carry_23_port, CO => 
                           position1_sub_216_I3_carry_24_port, S => 
                           position1_N1648);
   position1_sub_216_I4_U2_6 : ADD32 port map( A => position1_N1656, B => n37, 
                           CI => position1_sub_216_I4_carry_6_port, CO => 
                           position1_sub_216_I4_carry_7_port, S => 
                           position1_N1683);
   position1_sub_216_I4_U2_7 : ADD32 port map( A => position1_N1657, B => n67, 
                           CI => position1_sub_216_I4_carry_7_port, CO => 
                           position1_sub_216_I4_carry_8_port, S => 
                           position1_N1684);
   position1_sub_216_I4_U2_8 : ADD32 port map( A => position1_N1658, B => n38, 
                           CI => position1_sub_216_I4_carry_8_port, CO => 
                           position1_sub_216_I4_carry_9_port, S => 
                           position1_N1685);
   position1_sub_216_I4_U2_9 : ADD32 port map( A => position1_N1659, B => n276,
                           CI => position1_sub_216_I4_carry_9_port, CO => 
                           position1_sub_216_I4_carry_10_port, S => 
                           position1_N1686);
   position1_sub_216_I4_U2_10 : ADD32 port map( A => position1_N1660, B => n250
                           , CI => position1_sub_216_I4_carry_10_port, CO => 
                           position1_sub_216_I4_carry_11_port, S => 
                           position1_N1687);
   position1_sub_216_I4_U2_11 : ADD32 port map( A => position1_N1661, B => n280
                           , CI => position1_sub_216_I4_carry_11_port, CO => 
                           position1_sub_216_I4_carry_12_port, S => 
                           position1_N1688);
   position1_sub_216_I4_U2_12 : ADD32 port map( A => position1_N1662, B => n101
                           , CI => position1_sub_216_I4_carry_12_port, CO => 
                           position1_sub_216_I4_carry_13_port, S => 
                           position1_N1689);
   position1_sub_216_I4_U2_13 : ADD32 port map( A => position1_N1663, B => n256
                           , CI => position1_sub_216_I4_carry_13_port, CO => 
                           position1_sub_216_I4_carry_14_port, S => 
                           position1_N1690);
   position1_sub_216_I4_U2_14 : ADD32 port map( A => position1_N1664, B => n36,
                           CI => position1_sub_216_I4_carry_14_port, CO => 
                           position1_sub_216_I4_carry_15_port, S => 
                           position1_N1691);
   position1_sub_216_I4_U2_15 : ADD32 port map( A => position1_N1665, B => n288
                           , CI => position1_sub_216_I4_carry_15_port, CO => 
                           position1_sub_216_I4_carry_16_port, S => 
                           position1_N1692);
   position1_sub_216_I4_U2_16 : ADD32 port map( A => position1_N1666, B => n39,
                           CI => position1_sub_216_I4_carry_16_port, CO => 
                           position1_sub_216_I4_carry_17_port, S => 
                           position1_N1693);
   position1_sub_216_I4_U2_17 : ADD32 port map( A => position1_N1667, B => n263
                           , CI => position1_sub_216_I4_carry_17_port, CO => 
                           position1_sub_216_I4_carry_18_port, S => 
                           position1_N1694);
   position1_sub_216_I4_U2_18 : ADD32 port map( A => position1_N1668, B => n40,
                           CI => position1_sub_216_I4_carry_18_port, CO => 
                           position1_sub_216_I4_carry_19_port, S => 
                           position1_N1695);
   position1_sub_216_I4_U2_19 : ADD32 port map( A => position1_N1669, B => n296
                           , CI => position1_sub_216_I4_carry_19_port, CO => 
                           position1_sub_216_I4_carry_20_port, S => 
                           position1_N1696);
   position1_sub_216_I4_U2_20 : ADD32 port map( A => position1_N1670, B => n298
                           , CI => position1_sub_216_I4_carry_20_port, CO => 
                           position1_sub_216_I4_carry_21_port, S => 
                           position1_N1697);
   position1_sub_216_I4_U2_21 : ADD32 port map( A => position1_N1671, B => n300
                           , CI => position1_sub_216_I4_carry_21_port, CO => 
                           position1_sub_216_I4_carry_22_port, S => 
                           position1_N1698);
   position1_sub_216_I4_U2_22 : ADD32 port map( A => position1_N1672, B => n589
                           , CI => position1_sub_216_I4_carry_22_port, CO => 
                           position1_sub_216_I4_carry_23_port, S => 
                           position1_N1699);
   position1_sub_216_I5_U2_5 : ADD32 port map( A => n1239, B => n37, CI => 
                           position1_sub_216_I5_carry_5_port, CO => 
                           position1_sub_216_I5_carry_6_port, S => 
                           position1_N1734);
   position1_sub_216_I5_U2_6 : ADD32 port map( A => n1237, B => n245, CI => 
                           position1_sub_216_I5_carry_6_port, CO => 
                           position1_sub_216_I5_carry_7_port, S => 
                           position1_N1735);
   position1_sub_216_I5_U2_7 : ADD32 port map( A => n1235, B => n246, CI => 
                           position1_sub_216_I5_carry_7_port, CO => 
                           position1_sub_216_I5_carry_8_port, S => 
                           position1_N1736);
   position1_sub_216_I5_U2_8 : ADD32 port map( A => n1233, B => n248, CI => 
                           position1_sub_216_I5_carry_8_port, CO => 
                           position1_sub_216_I5_carry_9_port, S => 
                           position1_N1737);
   position1_sub_216_I5_U2_9 : ADD32 port map( A => n1231, B => n48, CI => 
                           position1_sub_216_I5_carry_9_port, CO => 
                           position1_sub_216_I5_carry_10_port, S => 
                           position1_N1738);
   position1_sub_216_I5_U2_10 : ADD32 port map( A => n1230, B => n252, CI => 
                           position1_sub_216_I5_carry_10_port, CO => 
                           position1_sub_216_I5_carry_11_port, S => 
                           position1_N1739);
   position1_sub_216_I5_U2_11 : ADD32 port map( A => n1228, B => n101, CI => 
                           position1_sub_216_I5_carry_11_port, CO => 
                           position1_sub_216_I5_carry_12_port, S => 
                           position1_N1740);
   position1_sub_216_I5_U2_12 : ADD32 port map( A => n1227, B => n284, CI => 
                           position1_sub_216_I5_carry_12_port, CO => 
                           position1_sub_216_I5_carry_13_port, S => 
                           position1_N1741);
   position1_sub_216_I5_U2_13 : ADD32 port map( A => n1226, B => n36, CI => 
                           position1_sub_216_I5_carry_13_port, CO => 
                           position1_sub_216_I5_carry_14_port, S => 
                           position1_N1742);
   position1_sub_216_I5_U2_14 : ADD32 port map( A => n1225, B => n259, CI => 
                           position1_sub_216_I5_carry_14_port, CO => 
                           position1_sub_216_I5_carry_15_port, S => 
                           position1_N1743);
   position1_sub_216_I5_U2_15 : ADD32 port map( A => n1224, B => n261, CI => 
                           position1_sub_216_I5_carry_15_port, CO => 
                           position1_sub_216_I5_carry_16_port, S => 
                           position1_N1744);
   position1_sub_216_I5_U2_16 : ADD32 port map( A => n1223, B => n292, CI => 
                           position1_sub_216_I5_carry_16_port, CO => 
                           position1_sub_216_I5_carry_17_port, S => 
                           position1_N1745);
   position1_sub_216_I5_U2_17 : ADD32 port map( A => n1222, B => n265, CI => 
                           position1_sub_216_I5_carry_17_port, CO => 
                           position1_sub_216_I5_carry_18_port, S => 
                           position1_N1746);
   position1_sub_216_I5_U2_18 : ADD32 port map( A => n1221, B => n267, CI => 
                           position1_sub_216_I5_carry_18_port, CO => 
                           position1_sub_216_I5_carry_19_port, S => 
                           position1_N1747);
   position1_sub_216_I5_U2_19 : ADD32 port map( A => n1220, B => n68, CI => 
                           position1_sub_216_I5_carry_19_port, CO => 
                           position1_sub_216_I5_carry_20_port, S => 
                           position1_N1748);
   position1_sub_216_I5_U2_20 : ADD32 port map( A => n1219, B => n45, CI => 
                           position1_sub_216_I5_carry_20_port, CO => 
                           position1_sub_216_I5_carry_21_port, S => 
                           position1_N1749);
   position1_sub_216_I5_U2_21 : ADD32 port map( A => n1218, B => n590, CI => 
                           position1_sub_216_I5_carry_21_port, CO => 
                           position1_sub_216_I5_carry_22_port, S => 
                           position1_N1750);
   position1_sub_216_I6_U2_4 : ADD32 port map( A => n1209, B => n37, CI => 
                           position1_sub_216_I6_carry_4_port, CO => 
                           position1_sub_216_I6_carry_5_port, S => 
                           position1_N1785);
   position1_sub_216_I6_U2_5 : ADD32 port map( A => n1208, B => n67, CI => 
                           position1_sub_216_I6_carry_5_port, CO => 
                           position1_sub_216_I6_carry_6_port, S => 
                           position1_N1786);
   position1_sub_216_I6_U2_6 : ADD32 port map( A => n1207, B => n38, CI => 
                           position1_sub_216_I6_carry_6_port, CO => 
                           position1_sub_216_I6_carry_7_port, S => 
                           position1_N1787);
   position1_sub_216_I6_U2_7 : ADD32 port map( A => n1206, B => n276, CI => 
                           position1_sub_216_I6_carry_7_port, CO => 
                           position1_sub_216_I6_carry_8_port, S => 
                           position1_N1788);
   position1_sub_216_I6_U2_8 : ADD32 port map( A => n1205, B => n48, CI => 
                           position1_sub_216_I6_carry_8_port, CO => 
                           position1_sub_216_I6_carry_9_port, S => 
                           position1_N1789);
   position1_sub_216_I6_U2_9 : ADD32 port map( A => n1204, B => n280, CI => 
                           position1_sub_216_I6_carry_9_port, CO => 
                           position1_sub_216_I6_carry_10_port, S => 
                           position1_N1790);
   position1_sub_216_I6_U2_10 : ADD32 port map( A => n1203, B => n101, CI => 
                           position1_sub_216_I6_carry_10_port, CO => 
                           position1_sub_216_I6_carry_11_port, S => 
                           position1_N1791);
   position1_sub_216_I6_U2_11 : ADD32 port map( A => n1202, B => n256, CI => 
                           position1_sub_216_I6_carry_11_port, CO => 
                           position1_sub_216_I6_carry_12_port, S => 
                           position1_N1792);
   position1_sub_216_I6_U2_12 : ADD32 port map( A => n1201, B => n36, CI => 
                           position1_sub_216_I6_carry_12_port, CO => 
                           position1_sub_216_I6_carry_13_port, S => 
                           position1_N1793);
   position1_sub_216_I6_U2_13 : ADD32 port map( A => n1200, B => n288, CI => 
                           position1_sub_216_I6_carry_13_port, CO => 
                           position1_sub_216_I6_carry_14_port, S => 
                           position1_N1794);
   position1_sub_216_I6_U2_14 : ADD32 port map( A => n1199, B => n39, CI => 
                           position1_sub_216_I6_carry_14_port, CO => 
                           position1_sub_216_I6_carry_15_port, S => 
                           position1_N1795);
   position1_sub_216_I6_U2_15 : ADD32 port map( A => n1198, B => n263, CI => 
                           position1_sub_216_I6_carry_15_port, CO => 
                           position1_sub_216_I6_carry_16_port, S => 
                           position1_N1796);
   position1_sub_216_I6_U2_16 : ADD32 port map( A => n1197, B => n40, CI => 
                           position1_sub_216_I6_carry_16_port, CO => 
                           position1_sub_216_I6_carry_17_port, S => 
                           position1_N1797);
   position1_sub_216_I6_U2_17 : ADD32 port map( A => n1196, B => n296, CI => 
                           position1_sub_216_I6_carry_17_port, CO => 
                           position1_sub_216_I6_carry_18_port, S => 
                           position1_N1798);
   position1_sub_216_I6_U2_18 : ADD32 port map( A => n1194, B => n68, CI => 
                           position1_sub_216_I6_carry_18_port, CO => 
                           position1_sub_216_I6_carry_19_port, S => 
                           position1_N1799);
   position1_sub_216_I6_U2_19 : ADD32 port map( A => n1193, B => n300, CI => 
                           position1_sub_216_I6_carry_19_port, CO => 
                           position1_sub_216_I6_carry_20_port, S => 
                           position1_N1800);
   position1_sub_216_I6_U2_20 : ADD32 port map( A => n1191, B => n590, CI => 
                           position1_sub_216_I6_carry_20_port, CO => 
                           position1_sub_216_I6_carry_21_port, S => 
                           position1_N1801);
   position1_sub_216_I7_U2_3 : ADD32 port map( A => n1182, B => n630, CI => 
                           position1_sub_216_I7_carry_3_port, CO => 
                           position1_sub_216_I7_carry_4_port, S => 
                           position1_N1836);
   position1_sub_216_I7_U2_4 : ADD32 port map( A => n1181, B => n67, CI => 
                           position1_sub_216_I7_carry_4_port, CO => 
                           position1_sub_216_I7_carry_5_port, S => 
                           position1_N1837);
   position1_sub_216_I7_U2_5 : ADD32 port map( A => n1180, B => n38, CI => 
                           position1_sub_216_I7_carry_5_port, CO => 
                           position1_sub_216_I7_carry_6_port, S => 
                           position1_N1838);
   position1_sub_216_I7_U2_6 : ADD32 port map( A => n1179, B => n248, CI => 
                           position1_sub_216_I7_carry_6_port, CO => 
                           position1_sub_216_I7_carry_7_port, S => 
                           position1_N1839);
   position1_sub_216_I7_U2_7 : ADD32 port map( A => n1178, B => n48, CI => 
                           position1_sub_216_I7_carry_7_port, CO => 
                           position1_sub_216_I7_carry_8_port, S => 
                           position1_N1840);
   position1_sub_216_I7_U2_8 : ADD32 port map( A => n1177, B => n252, CI => 
                           position1_sub_216_I7_carry_8_port, CO => 
                           position1_sub_216_I7_carry_9_port, S => 
                           position1_N1841);
   position1_sub_216_I7_U2_9 : ADD32 port map( A => n1176, B => n101, CI => 
                           position1_sub_216_I7_carry_9_port, CO => 
                           position1_sub_216_I7_carry_10_port, S => 
                           position1_N1842);
   position1_sub_216_I7_U2_10 : ADD32 port map( A => n1175, B => n284, CI => 
                           position1_sub_216_I7_carry_10_port, CO => 
                           position1_sub_216_I7_carry_11_port, S => 
                           position1_N1843);
   position1_sub_216_I7_U2_11 : ADD32 port map( A => n1174, B => n36, CI => 
                           position1_sub_216_I7_carry_11_port, CO => 
                           position1_sub_216_I7_carry_12_port, S => 
                           position1_N1844);
   position1_sub_216_I7_U2_12 : ADD32 port map( A => n1173, B => n259, CI => 
                           position1_sub_216_I7_carry_12_port, CO => 
                           position1_sub_216_I7_carry_13_port, S => 
                           position1_N1845);
   position1_sub_216_I7_U2_13 : ADD32 port map( A => n1172, B => n39, CI => 
                           position1_sub_216_I7_carry_13_port, CO => 
                           position1_sub_216_I7_carry_14_port, S => 
                           position1_N1846);
   position1_sub_216_I7_U2_14 : ADD32 port map( A => n1171, B => n292, CI => 
                           position1_sub_216_I7_carry_14_port, CO => 
                           position1_sub_216_I7_carry_15_port, S => 
                           position1_N1847);
   position1_sub_216_I7_U2_15 : ADD32 port map( A => n1170, B => n40, CI => 
                           position1_sub_216_I7_carry_15_port, CO => 
                           position1_sub_216_I7_carry_16_port, S => 
                           position1_N1848);
   position1_sub_216_I7_U2_16 : ADD32 port map( A => n1169, B => n296, CI => 
                           position1_sub_216_I7_carry_16_port, CO => 
                           position1_sub_216_I7_carry_17_port, S => 
                           position1_N1849);
   position1_sub_216_I7_U2_17 : ADD32 port map( A => n1168, B => n68, CI => 
                           position1_sub_216_I7_carry_17_port, CO => 
                           position1_sub_216_I7_carry_18_port, S => 
                           position1_N1850);
   position1_sub_216_I7_U2_18 : ADD32 port map( A => n1167, B => n45, CI => 
                           position1_sub_216_I7_carry_18_port, CO => 
                           position1_sub_216_I7_carry_19_port, S => 
                           position1_N1851);
   position1_sub_216_I7_U2_19 : ADD32 port map( A => n1166, B => n590, CI => 
                           position1_sub_216_I7_carry_19_port, CO => 
                           position1_sub_216_I7_carry_20_port, S => 
                           position1_N1852);
   position1_sub_216_I8_U2_2 : ADD32 port map( A => n1157, B => n37, CI => 
                           position1_sub_216_I8_carry_2_port, CO => 
                           position1_sub_216_I8_carry_3_port, S => 
                           position1_N1887);
   position1_sub_216_I8_U2_3 : ADD32 port map( A => n1155, B => n67, CI => 
                           position1_sub_216_I8_carry_3_port, CO => 
                           position1_sub_216_I8_carry_4_port, S => 
                           position1_N1888);
   position1_sub_216_I8_U2_4 : ADD32 port map( A => n1154, B => n38, CI => 
                           position1_sub_216_I8_carry_4_port, CO => 
                           position1_sub_216_I8_carry_5_port, S => 
                           position1_N1889);
   position1_sub_216_I8_U2_5 : ADD32 port map( A => n1152, B => n276, CI => 
                           position1_sub_216_I8_carry_5_port, CO => 
                           position1_sub_216_I8_carry_6_port, S => 
                           position1_N1890);
   position1_sub_216_I8_U2_6 : ADD32 port map( A => n1151, B => n48, CI => 
                           position1_sub_216_I8_carry_6_port, CO => 
                           position1_sub_216_I8_carry_7_port, S => 
                           position1_N1891);
   position1_sub_216_I8_U2_7 : ADD32 port map( A => n1149, B => n280, CI => 
                           position1_sub_216_I8_carry_7_port, CO => 
                           position1_sub_216_I8_carry_8_port, S => 
                           position1_N1892);
   position1_sub_216_I8_U2_8 : ADD32 port map( A => n1148, B => n101, CI => 
                           position1_sub_216_I8_carry_8_port, CO => 
                           position1_sub_216_I8_carry_9_port, S => 
                           position1_N1893);
   position1_sub_216_I8_U2_9 : ADD32 port map( A => n1146, B => n284, CI => 
                           position1_sub_216_I8_carry_9_port, CO => 
                           position1_sub_216_I8_carry_10_port, S => 
                           position1_N1894);
   position1_sub_216_I8_U2_10 : ADD32 port map( A => n1145, B => n36, CI => 
                           position1_sub_216_I8_carry_10_port, CO => 
                           position1_sub_216_I8_carry_11_port, S => 
                           position1_N1895);
   position1_sub_216_I8_U2_11 : ADD32 port map( A => n1144, B => n288, CI => 
                           position1_sub_216_I8_carry_11_port, CO => 
                           position1_sub_216_I8_carry_12_port, S => 
                           position1_N1896);
   position1_sub_216_I8_U2_12 : ADD32 port map( A => n1142, B => n39, CI => 
                           position1_sub_216_I8_carry_12_port, CO => 
                           position1_sub_216_I8_carry_13_port, S => 
                           position1_N1897);
   position1_sub_216_I8_U2_13 : ADD32 port map( A => n1140, B => n292, CI => 
                           position1_sub_216_I8_carry_13_port, CO => 
                           position1_sub_216_I8_carry_14_port, S => 
                           position1_N1898);
   position1_sub_216_I8_U2_14 : ADD32 port map( A => n1139, B => n40, CI => 
                           position1_sub_216_I8_carry_14_port, CO => 
                           position1_sub_216_I8_carry_15_port, S => 
                           position1_N1899);
   position1_sub_216_I8_U2_15 : ADD32 port map( A => n1137, B => n296, CI => 
                           position1_sub_216_I8_carry_15_port, CO => 
                           position1_sub_216_I8_carry_16_port, S => 
                           position1_N1900);
   position1_sub_216_I8_U2_16 : ADD32 port map( A => n1136, B => n68, CI => 
                           position1_sub_216_I8_carry_16_port, CO => 
                           position1_sub_216_I8_carry_17_port, S => 
                           position1_N1901);
   position1_sub_216_I8_U2_17 : ADD32 port map( A => n1135, B => n45, CI => 
                           position1_sub_216_I8_carry_17_port, CO => 
                           position1_sub_216_I8_carry_18_port, S => 
                           position1_N1902);
   position1_sub_216_I8_U2_18 : ADD32 port map( A => n1134, B => n590, CI => 
                           position1_sub_216_I8_carry_18_port, CO => 
                           position1_sub_216_I8_carry_19_port, S => 
                           position1_N1903);
   position1_sub_226_U2_9 : ADD32 port map( A => position1_y_sum_9_port, B => 
                           n37, CI => position1_sub_226_carry_9_port, CO => 
                           position1_sub_226_carry_10_port, S => 
                           position1_N1947);
   position1_sub_226_U2_10 : ADD32 port map( A => position1_y_sum_10_port, B =>
                           n67, CI => position1_sub_226_carry_10_port, CO => 
                           position1_sub_226_carry_11_port, S => 
                           position1_N1948);
   position1_sub_226_U2_11 : ADD32 port map( A => position1_y_sum_11_port, B =>
                           n38, CI => position1_sub_226_carry_11_port, CO => 
                           position1_sub_226_carry_12_port, S => 
                           position1_N1949);
   position1_sub_226_U2_12 : ADD32 port map( A => position1_y_sum_12_port, B =>
                           n42, CI => position1_sub_226_carry_12_port, CO => 
                           position1_sub_226_carry_13_port, S => 
                           position1_N1950);
   position1_sub_226_U2_13 : ADD32 port map( A => position1_y_sum_13_port, B =>
                           n48, CI => position1_sub_226_carry_13_port, CO => 
                           position1_sub_226_carry_14_port, S => 
                           position1_N1951);
   position1_sub_226_U2_14 : ADD32 port map( A => position1_y_sum_14_port, B =>
                           n46, CI => position1_sub_226_carry_14_port, CO => 
                           position1_sub_226_carry_15_port, S => 
                           position1_N1952);
   position1_sub_226_U2_15 : ADD32 port map( A => position1_y_sum_15_port, B =>
                           n101, CI => position1_sub_226_carry_15_port, CO => 
                           position1_sub_226_carry_16_port, S => 
                           position1_N1953);
   position1_sub_226_U2_16 : ADD32 port map( A => position1_y_sum_16_port, B =>
                           n41, CI => position1_sub_226_carry_16_port, CO => 
                           position1_sub_226_carry_17_port, S => 
                           position1_N1954);
   position1_sub_226_U2_17 : ADD32 port map( A => position1_y_sum_17_port, B =>
                           n36, CI => position1_sub_226_carry_17_port, CO => 
                           position1_sub_226_carry_18_port, S => 
                           position1_N1955);
   position1_sub_226_U2_18 : ADD32 port map( A => position1_y_sum_18_port, B =>
                           n288, CI => position1_sub_226_carry_18_port, CO => 
                           position1_sub_226_carry_19_port, S => 
                           position1_N1956);
   position1_sub_226_U2_19 : ADD32 port map( A => position1_y_sum_19_port, B =>
                           n39, CI => position1_sub_226_carry_19_port, CO => 
                           position1_sub_226_carry_20_port, S => 
                           position1_N1957);
   position1_sub_226_U2_20 : ADD32 port map( A => position1_y_sum_20_port, B =>
                           n44, CI => position1_sub_226_carry_20_port, CO => 
                           position1_sub_226_carry_21_port, S => 
                           position1_N1958);
   position1_sub_226_U2_21 : ADD32 port map( A => position1_y_sum_21_port, B =>
                           n40, CI => position1_sub_226_carry_21_port, CO => 
                           position1_sub_226_carry_22_port, S => 
                           position1_N1959);
   position1_sub_226_U2_22 : ADD32 port map( A => position1_y_sum_22_port, B =>
                           n43, CI => position1_sub_226_carry_22_port, CO => 
                           position1_sub_226_carry_23_port, S => 
                           position1_N1960);
   position1_sub_226_U2_23 : ADD32 port map( A => position1_y_sum_23_port, B =>
                           n68, CI => position1_sub_226_carry_23_port, CO => 
                           position1_sub_226_carry_24_port, S => 
                           position1_N1961);
   position1_sub_226_I2_U2_8 : ADD32 port map( A => position1_N1971, B => n630,
                           CI => position1_sub_226_I2_carry_8_port, CO => 
                           position1_sub_226_I2_carry_9_port, S => 
                           position1_N1998);
   position1_sub_226_I2_U2_9 : ADD32 port map( A => position1_N1972, B => n67, 
                           CI => position1_sub_226_I2_carry_9_port, CO => 
                           position1_sub_226_I2_carry_10_port, S => 
                           position1_N1999);
   position1_sub_226_I2_U2_10 : ADD32 port map( A => position1_N1973, B => n38,
                           CI => position1_sub_226_I2_carry_10_port, CO => 
                           position1_sub_226_I2_carry_11_port, S => 
                           position1_N2000);
   position1_sub_226_I2_U2_11 : ADD32 port map( A => position1_N1974, B => n42,
                           CI => position1_sub_226_I2_carry_11_port, CO => 
                           position1_sub_226_I2_carry_12_port, S => 
                           position1_N2001);
   position1_sub_226_I2_U2_12 : ADD32 port map( A => position1_N1975, B => n48,
                           CI => position1_sub_226_I2_carry_12_port, CO => 
                           position1_sub_226_I2_carry_13_port, S => 
                           position1_N2002);
   position1_sub_226_I2_U2_13 : ADD32 port map( A => position1_N1976, B => n46,
                           CI => position1_sub_226_I2_carry_13_port, CO => 
                           position1_sub_226_I2_carry_14_port, S => 
                           position1_N2003);
   position1_sub_226_I2_U2_14 : ADD32 port map( A => position1_N1977, B => n101
                           , CI => position1_sub_226_I2_carry_14_port, CO => 
                           position1_sub_226_I2_carry_15_port, S => 
                           position1_N2004);
   position1_sub_226_I2_U2_15 : ADD32 port map( A => position1_N1978, B => n41,
                           CI => position1_sub_226_I2_carry_15_port, CO => 
                           position1_sub_226_I2_carry_16_port, S => 
                           position1_N2005);
   position1_sub_226_I2_U2_16 : ADD32 port map( A => position1_N1979, B => n36,
                           CI => position1_sub_226_I2_carry_16_port, CO => 
                           position1_sub_226_I2_carry_17_port, S => 
                           position1_N2006);
   position1_sub_226_I2_U2_17 : ADD32 port map( A => position1_N1980, B => n47,
                           CI => position1_sub_226_I2_carry_17_port, CO => 
                           position1_sub_226_I2_carry_18_port, S => 
                           position1_N2007);
   position1_sub_226_I2_U2_18 : ADD32 port map( A => position1_N1981, B => n39,
                           CI => position1_sub_226_I2_carry_18_port, CO => 
                           position1_sub_226_I2_carry_19_port, S => 
                           position1_N2008);
   position1_sub_226_I2_U2_19 : ADD32 port map( A => position1_N1982, B => n44,
                           CI => position1_sub_226_I2_carry_19_port, CO => 
                           position1_sub_226_I2_carry_20_port, S => 
                           position1_N2009);
   position1_sub_226_I2_U2_20 : ADD32 port map( A => position1_N1983, B => n40,
                           CI => position1_sub_226_I2_carry_20_port, CO => 
                           position1_sub_226_I2_carry_21_port, S => 
                           position1_N2010);
   position1_sub_226_I2_U2_21 : ADD32 port map( A => position1_N1984, B => n43,
                           CI => position1_sub_226_I2_carry_21_port, CO => 
                           position1_sub_226_I2_carry_22_port, S => 
                           position1_N2011);
   position1_sub_226_I2_U2_22 : ADD32 port map( A => position1_N1985, B => n68,
                           CI => position1_sub_226_I2_carry_22_port, CO => 
                           position1_sub_226_I2_carry_23_port, S => 
                           position1_N2012);
   position1_sub_226_I2_U2_23 : ADD32 port map( A => position1_N1986, B => n45,
                           CI => position1_sub_226_I2_carry_23_port, CO => 
                           position1_sub_226_I2_carry_24_port, S => 
                           position1_N2013);
   position1_sub_226_I3_U2_7 : ADD32 port map( A => n1081, B => n37, CI => 
                           position1_sub_226_I3_carry_7_port, CO => 
                           position1_sub_226_I3_carry_8_port, S => 
                           position1_N2049);
   position1_sub_226_I3_U2_8 : ADD32 port map( A => n1079, B => n67, CI => 
                           position1_sub_226_I3_carry_8_port, CO => 
                           position1_sub_226_I3_carry_9_port, S => 
                           position1_N2050);
   position1_sub_226_I3_U2_9 : ADD32 port map( A => n1076, B => n38, CI => 
                           position1_sub_226_I3_carry_9_port, CO => 
                           position1_sub_226_I3_carry_10_port, S => 
                           position1_N2051);
   position1_sub_226_I3_U2_10 : ADD32 port map( A => n1074, B => n42, CI => 
                           position1_sub_226_I3_carry_10_port, CO => 
                           position1_sub_226_I3_carry_11_port, S => 
                           position1_N2052);
   position1_sub_226_I3_U2_11 : ADD32 port map( A => n1071, B => n48, CI => 
                           position1_sub_226_I3_carry_11_port, CO => 
                           position1_sub_226_I3_carry_12_port, S => 
                           position1_N2053);
   position1_sub_226_I3_U2_12 : ADD32 port map( A => n1069, B => n46, CI => 
                           position1_sub_226_I3_carry_12_port, CO => 
                           position1_sub_226_I3_carry_13_port, S => 
                           position1_N2054);
   position1_sub_226_I3_U2_13 : ADD32 port map( A => n1067, B => n101, CI => 
                           position1_sub_226_I3_carry_13_port, CO => 
                           position1_sub_226_I3_carry_14_port, S => 
                           position1_N2055);
   position1_sub_226_I3_U2_14 : ADD32 port map( A => n1065, B => n41, CI => 
                           position1_sub_226_I3_carry_14_port, CO => 
                           position1_sub_226_I3_carry_15_port, S => 
                           position1_N2056);
   position1_sub_226_I3_U2_15 : ADD32 port map( A => n1063, B => n36, CI => 
                           position1_sub_226_I3_carry_15_port, CO => 
                           position1_sub_226_I3_carry_16_port, S => 
                           position1_N2057);
   position1_sub_226_I3_U2_16 : ADD32 port map( A => n1061, B => n47, CI => 
                           position1_sub_226_I3_carry_16_port, CO => 
                           position1_sub_226_I3_carry_17_port, S => 
                           position1_N2058);
   position1_sub_226_I3_U2_17 : ADD32 port map( A => n1059, B => n39, CI => 
                           position1_sub_226_I3_carry_17_port, CO => 
                           position1_sub_226_I3_carry_18_port, S => 
                           position1_N2059);
   position1_sub_226_I3_U2_18 : ADD32 port map( A => n1057, B => n44, CI => 
                           position1_sub_226_I3_carry_18_port, CO => 
                           position1_sub_226_I3_carry_19_port, S => 
                           position1_N2060);
   position1_sub_226_I3_U2_19 : ADD32 port map( A => n1055, B => n40, CI => 
                           position1_sub_226_I3_carry_19_port, CO => 
                           position1_sub_226_I3_carry_20_port, S => 
                           position1_N2061);
   position1_sub_226_I3_U2_20 : ADD32 port map( A => n1053, B => n43, CI => 
                           position1_sub_226_I3_carry_20_port, CO => 
                           position1_sub_226_I3_carry_21_port, S => 
                           position1_N2062);
   position1_sub_226_I3_U2_21 : ADD32 port map( A => n1051, B => n68, CI => 
                           position1_sub_226_I3_carry_21_port, CO => 
                           position1_sub_226_I3_carry_22_port, S => 
                           position1_N2063);
   position1_sub_226_I3_U2_22 : ADD32 port map( A => n1050, B => n45, CI => 
                           position1_sub_226_I3_carry_22_port, CO => 
                           position1_sub_226_I3_carry_23_port, S => 
                           position1_N2064);
   position1_sub_226_I3_U2_23 : ADD32 port map( A => n1049, B => n591, CI => 
                           position1_sub_226_I3_carry_23_port, CO => 
                           position1_sub_226_I3_carry_24_port, S => 
                           position1_N2065);
   position1_sub_226_I4_U2_6 : ADD32 port map( A => position1_N2073, B => n630,
                           CI => position1_sub_226_I4_carry_6_port, CO => 
                           position1_sub_226_I4_carry_7_port, S => 
                           position1_N2100);
   position1_sub_226_I4_U2_7 : ADD32 port map( A => position1_N2074, B => n67, 
                           CI => position1_sub_226_I4_carry_7_port, CO => 
                           position1_sub_226_I4_carry_8_port, S => 
                           position1_N2101);
   position1_sub_226_I4_U2_8 : ADD32 port map( A => position1_N2075, B => n38, 
                           CI => position1_sub_226_I4_carry_8_port, CO => 
                           position1_sub_226_I4_carry_9_port, S => 
                           position1_N2102);
   position1_sub_226_I4_U2_9 : ADD32 port map( A => position1_N2076, B => n42, 
                           CI => position1_sub_226_I4_carry_9_port, CO => 
                           position1_sub_226_I4_carry_10_port, S => 
                           position1_N2103);
   position1_sub_226_I4_U2_10 : ADD32 port map( A => position1_N2077, B => n48,
                           CI => position1_sub_226_I4_carry_10_port, CO => 
                           position1_sub_226_I4_carry_11_port, S => 
                           position1_N2104);
   position1_sub_226_I4_U2_11 : ADD32 port map( A => position1_N2078, B => n46,
                           CI => position1_sub_226_I4_carry_11_port, CO => 
                           position1_sub_226_I4_carry_12_port, S => 
                           position1_N2105);
   position1_sub_226_I4_U2_12 : ADD32 port map( A => position1_N2079, B => n101
                           , CI => position1_sub_226_I4_carry_12_port, CO => 
                           position1_sub_226_I4_carry_13_port, S => 
                           position1_N2106);
   position1_sub_226_I4_U2_13 : ADD32 port map( A => position1_N2080, B => n41,
                           CI => position1_sub_226_I4_carry_13_port, CO => 
                           position1_sub_226_I4_carry_14_port, S => 
                           position1_N2107);
   position1_sub_226_I4_U2_14 : ADD32 port map( A => position1_N2081, B => n36,
                           CI => position1_sub_226_I4_carry_14_port, CO => 
                           position1_sub_226_I4_carry_15_port, S => 
                           position1_N2108);
   position1_sub_226_I4_U2_15 : ADD32 port map( A => position1_N2082, B => n47,
                           CI => position1_sub_226_I4_carry_15_port, CO => 
                           position1_sub_226_I4_carry_16_port, S => 
                           position1_N2109);
   position1_sub_226_I4_U2_16 : ADD32 port map( A => position1_N2083, B => n39,
                           CI => position1_sub_226_I4_carry_16_port, CO => 
                           position1_sub_226_I4_carry_17_port, S => 
                           position1_N2110);
   position1_sub_226_I4_U2_17 : ADD32 port map( A => position1_N2084, B => n44,
                           CI => position1_sub_226_I4_carry_17_port, CO => 
                           position1_sub_226_I4_carry_18_port, S => 
                           position1_N2111);
   position1_sub_226_I4_U2_18 : ADD32 port map( A => position1_N2085, B => n40,
                           CI => position1_sub_226_I4_carry_18_port, CO => 
                           position1_sub_226_I4_carry_19_port, S => 
                           position1_N2112);
   position1_sub_226_I4_U2_19 : ADD32 port map( A => position1_N2086, B => n43,
                           CI => position1_sub_226_I4_carry_19_port, CO => 
                           position1_sub_226_I4_carry_20_port, S => 
                           position1_N2113);
   position1_sub_226_I4_U2_20 : ADD32 port map( A => position1_N2087, B => n68,
                           CI => position1_sub_226_I4_carry_20_port, CO => 
                           position1_sub_226_I4_carry_21_port, S => 
                           position1_N2114);
   position1_sub_226_I4_U2_21 : ADD32 port map( A => position1_N2088, B => n45,
                           CI => position1_sub_226_I4_carry_21_port, CO => 
                           position1_sub_226_I4_carry_22_port, S => 
                           position1_N2115);
   position1_sub_226_I4_U2_22 : ADD32 port map( A => position1_N2089, B => n591
                           , CI => position1_sub_226_I4_carry_22_port, CO => 
                           position1_sub_226_I4_carry_23_port, S => 
                           position1_N2116);
   position1_sub_226_I5_U2_5 : ADD32 port map( A => n1020, B => n37, CI => 
                           position1_sub_226_I5_carry_5_port, CO => 
                           position1_sub_226_I5_carry_6_port, S => 
                           position1_N2151);
   position1_sub_226_I5_U2_6 : ADD32 port map( A => n1018, B => n245, CI => 
                           position1_sub_226_I5_carry_6_port, CO => 
                           position1_sub_226_I5_carry_7_port, S => 
                           position1_N2152);
   position1_sub_226_I5_U2_7 : ADD32 port map( A => n1016, B => n274, CI => 
                           position1_sub_226_I5_carry_7_port, CO => 
                           position1_sub_226_I5_carry_8_port, S => 
                           position1_N2153);
   position1_sub_226_I5_U2_8 : ADD32 port map( A => n1014, B => n42, CI => 
                           position1_sub_226_I5_carry_8_port, CO => 
                           position1_sub_226_I5_carry_9_port, S => 
                           position1_N2154);
   position1_sub_226_I5_U2_9 : ADD32 port map( A => n1012, B => n278, CI => 
                           position1_sub_226_I5_carry_9_port, CO => 
                           position1_sub_226_I5_carry_10_port, S => 
                           position1_N2155);
   position1_sub_226_I5_U2_10 : ADD32 port map( A => n1011, B => n46, CI => 
                           position1_sub_226_I5_carry_10_port, CO => 
                           position1_sub_226_I5_carry_11_port, S => 
                           position1_N2156);
   position1_sub_226_I5_U2_11 : ADD32 port map( A => n1009, B => n101, CI => 
                           position1_sub_226_I5_carry_11_port, CO => 
                           position1_sub_226_I5_carry_12_port, S => 
                           position1_N2157);
   position1_sub_226_I5_U2_12 : ADD32 port map( A => n1008, B => n41, CI => 
                           position1_sub_226_I5_carry_12_port, CO => 
                           position1_sub_226_I5_carry_13_port, S => 
                           position1_N2158);
   position1_sub_226_I5_U2_13 : ADD32 port map( A => n1007, B => n36, CI => 
                           position1_sub_226_I5_carry_13_port, CO => 
                           position1_sub_226_I5_carry_14_port, S => 
                           position1_N2159);
   position1_sub_226_I5_U2_14 : ADD32 port map( A => n1006, B => n47, CI => 
                           position1_sub_226_I5_carry_14_port, CO => 
                           position1_sub_226_I5_carry_15_port, S => 
                           position1_N2160);
   position1_sub_226_I5_U2_15 : ADD32 port map( A => n1005, B => n261, CI => 
                           position1_sub_226_I5_carry_15_port, CO => 
                           position1_sub_226_I5_carry_16_port, S => 
                           position1_N2161);
   position1_sub_226_I5_U2_16 : ADD32 port map( A => n1004, B => n292, CI => 
                           position1_sub_226_I5_carry_16_port, CO => 
                           position1_sub_226_I5_carry_17_port, S => 
                           position1_N2162);
   position1_sub_226_I5_U2_17 : ADD32 port map( A => n1003, B => n265, CI => 
                           position1_sub_226_I5_carry_17_port, CO => 
                           position1_sub_226_I5_carry_18_port, S => 
                           position1_N2163);
   position1_sub_226_I5_U2_18 : ADD32 port map( A => n1002, B => n267, CI => 
                           position1_sub_226_I5_carry_18_port, CO => 
                           position1_sub_226_I5_carry_19_port, S => 
                           position1_N2164);
   position1_sub_226_I5_U2_19 : ADD32 port map( A => n1001, B => n269, CI => 
                           position1_sub_226_I5_carry_19_port, CO => 
                           position1_sub_226_I5_carry_20_port, S => 
                           position1_N2165);
   position1_sub_226_I5_U2_20 : ADD32 port map( A => n1000, B => n300, CI => 
                           position1_sub_226_I5_carry_20_port, CO => 
                           position1_sub_226_I5_carry_21_port, S => 
                           position1_N2166);
   position1_sub_226_I5_U2_21 : ADD32 port map( A => n999, B => n591, CI => 
                           position1_sub_226_I5_carry_21_port, CO => 
                           position1_sub_226_I5_carry_22_port, S => 
                           position1_N2167);
   position1_sub_226_I6_U2_4 : ADD32 port map( A => n990, B => n37, CI => 
                           position1_sub_226_I6_carry_4_port, CO => 
                           position1_sub_226_I6_carry_5_port, S => 
                           position1_N2202);
   position1_sub_226_I6_U2_5 : ADD32 port map( A => n989, B => n272, CI => 
                           position1_sub_226_I6_carry_5_port, CO => 
                           position1_sub_226_I6_carry_6_port, S => 
                           position1_N2203);
   position1_sub_226_I6_U2_6 : ADD32 port map( A => n988, B => n246, CI => 
                           position1_sub_226_I6_carry_6_port, CO => 
                           position1_sub_226_I6_carry_7_port, S => 
                           position1_N2204);
   position1_sub_226_I6_U2_7 : ADD32 port map( A => n987, B => n42, CI => 
                           position1_sub_226_I6_carry_7_port, CO => 
                           position1_sub_226_I6_carry_8_port, S => 
                           position1_N2205);
   position1_sub_226_I6_U2_8 : ADD32 port map( A => n986, B => n250, CI => 
                           position1_sub_226_I6_carry_8_port, CO => 
                           position1_sub_226_I6_carry_9_port, S => 
                           position1_N2206);
   position1_sub_226_I6_U2_9 : ADD32 port map( A => n985, B => n46, CI => 
                           position1_sub_226_I6_carry_9_port, CO => 
                           position1_sub_226_I6_carry_10_port, S => 
                           position1_N2207);
   position1_sub_226_I6_U2_10 : ADD32 port map( A => n984, B => n254, CI => 
                           position1_sub_226_I6_carry_10_port, CO => 
                           position1_sub_226_I6_carry_11_port, S => 
                           position1_N2208);
   position1_sub_226_I6_U2_11 : ADD32 port map( A => n983, B => n41, CI => 
                           position1_sub_226_I6_carry_11_port, CO => 
                           position1_sub_226_I6_carry_12_port, S => 
                           position1_N2209);
   position1_sub_226_I6_U2_12 : ADD32 port map( A => n982, B => n286, CI => 
                           position1_sub_226_I6_carry_12_port, CO => 
                           position1_sub_226_I6_carry_13_port, S => 
                           position1_N2210);
   position1_sub_226_I6_U2_13 : ADD32 port map( A => n981, B => n47, CI => 
                           position1_sub_226_I6_carry_13_port, CO => 
                           position1_sub_226_I6_carry_14_port, S => 
                           position1_N2211);
   position1_sub_226_I6_U2_14 : ADD32 port map( A => n980, B => n290, CI => 
                           position1_sub_226_I6_carry_14_port, CO => 
                           position1_sub_226_I6_carry_15_port, S => 
                           position1_N2212);
   position1_sub_226_I6_U2_15 : ADD32 port map( A => n979, B => n44, CI => 
                           position1_sub_226_I6_carry_15_port, CO => 
                           position1_sub_226_I6_carry_16_port, S => 
                           position1_N2213);
   position1_sub_226_I6_U2_16 : ADD32 port map( A => n978, B => n294, CI => 
                           position1_sub_226_I6_carry_16_port, CO => 
                           position1_sub_226_I6_carry_17_port, S => 
                           position1_N2214);
   position1_sub_226_I6_U2_17 : ADD32 port map( A => n977, B => n43, CI => 
                           position1_sub_226_I6_carry_17_port, CO => 
                           position1_sub_226_I6_carry_18_port, S => 
                           position1_N2215);
   position1_sub_226_I6_U2_18 : ADD32 port map( A => n975, B => n298, CI => 
                           position1_sub_226_I6_carry_18_port, CO => 
                           position1_sub_226_I6_carry_19_port, S => 
                           position1_N2216);
   position1_sub_226_I6_U2_19 : ADD32 port map( A => n974, B => n300, CI => 
                           position1_sub_226_I6_carry_19_port, CO => 
                           position1_sub_226_I6_carry_20_port, S => 
                           position1_N2217);
   position1_sub_226_I6_U2_20 : ADD32 port map( A => n972, B => n591, CI => 
                           position1_sub_226_I6_carry_20_port, CO => 
                           position1_sub_226_I6_carry_21_port, S => 
                           position1_N2218);
   position1_sub_226_I7_U2_3 : ADD32 port map( A => n963, B => n37, CI => 
                           position1_sub_226_I7_carry_3_port, CO => 
                           position1_sub_226_I7_carry_4_port, S => 
                           position1_N2253);
   position1_sub_226_I7_U2_4 : ADD32 port map( A => n962, B => n245, CI => 
                           position1_sub_226_I7_carry_4_port, CO => 
                           position1_sub_226_I7_carry_5_port, S => 
                           position1_N2254);
   position1_sub_226_I7_U2_5 : ADD32 port map( A => n961, B => n274, CI => 
                           position1_sub_226_I7_carry_5_port, CO => 
                           position1_sub_226_I7_carry_6_port, S => 
                           position1_N2255);
   position1_sub_226_I7_U2_6 : ADD32 port map( A => n960, B => n42, CI => 
                           position1_sub_226_I7_carry_6_port, CO => 
                           position1_sub_226_I7_carry_7_port, S => 
                           position1_N2256);
   position1_sub_226_I7_U2_7 : ADD32 port map( A => n959, B => n278, CI => 
                           position1_sub_226_I7_carry_7_port, CO => 
                           position1_sub_226_I7_carry_8_port, S => 
                           position1_N2257);
   position1_sub_226_I7_U2_8 : ADD32 port map( A => n958, B => n46, CI => 
                           position1_sub_226_I7_carry_8_port, CO => 
                           position1_sub_226_I7_carry_9_port, S => 
                           position1_N2258);
   position1_sub_226_I7_U2_9 : ADD32 port map( A => n957, B => n282, CI => 
                           position1_sub_226_I7_carry_9_port, CO => 
                           position1_sub_226_I7_carry_10_port, S => 
                           position1_N2259);
   position1_sub_226_I7_U2_10 : ADD32 port map( A => n956, B => n41, CI => 
                           position1_sub_226_I7_carry_10_port, CO => 
                           position1_sub_226_I7_carry_11_port, S => 
                           position1_N2260);
   position1_sub_226_I7_U2_11 : ADD32 port map( A => n955, B => n286, CI => 
                           position1_sub_226_I7_carry_11_port, CO => 
                           position1_sub_226_I7_carry_12_port, S => 
                           position1_N2261);
   position1_sub_226_I7_U2_12 : ADD32 port map( A => n954, B => n47, CI => 
                           position1_sub_226_I7_carry_12_port, CO => 
                           position1_sub_226_I7_carry_13_port, S => 
                           position1_N2262);
   position1_sub_226_I7_U2_13 : ADD32 port map( A => n953, B => n261, CI => 
                           position1_sub_226_I7_carry_13_port, CO => 
                           position1_sub_226_I7_carry_14_port, S => 
                           position1_N2263);
   position1_sub_226_I7_U2_14 : ADD32 port map( A => n952, B => n44, CI => 
                           position1_sub_226_I7_carry_14_port, CO => 
                           position1_sub_226_I7_carry_15_port, S => 
                           position1_N2264);
   position1_sub_226_I7_U2_15 : ADD32 port map( A => n951, B => n265, CI => 
                           position1_sub_226_I7_carry_15_port, CO => 
                           position1_sub_226_I7_carry_16_port, S => 
                           position1_N2265);
   position1_sub_226_I7_U2_16 : ADD32 port map( A => n950, B => n43, CI => 
                           position1_sub_226_I7_carry_16_port, CO => 
                           position1_sub_226_I7_carry_17_port, S => 
                           position1_N2266);
   position1_sub_226_I7_U2_17 : ADD32 port map( A => n949, B => n269, CI => 
                           position1_sub_226_I7_carry_17_port, CO => 
                           position1_sub_226_I7_carry_18_port, S => 
                           position1_N2267);
   position1_sub_226_I7_U2_18 : ADD32 port map( A => n948, B => n300, CI => 
                           position1_sub_226_I7_carry_18_port, CO => 
                           position1_sub_226_I7_carry_19_port, S => 
                           position1_N2268);
   position1_sub_226_I7_U2_19 : ADD32 port map( A => n947, B => n592, CI => 
                           position1_sub_226_I7_carry_19_port, CO => 
                           position1_sub_226_I7_carry_20_port, S => 
                           position1_N2269);
   position1_sub_226_I8_U2_2 : ADD32 port map( A => n938, B => n630, CI => 
                           position1_sub_226_I8_carry_2_port, CO => 
                           position1_sub_226_I8_carry_3_port, S => 
                           position1_N2304);
   position1_sub_226_I8_U2_3 : ADD32 port map( A => n936, B => n272, CI => 
                           position1_sub_226_I8_carry_3_port, CO => 
                           position1_sub_226_I8_carry_4_port, S => 
                           position1_N2305);
   position1_sub_226_I8_U2_4 : ADD32 port map( A => n935, B => n246, CI => 
                           position1_sub_226_I8_carry_4_port, CO => 
                           position1_sub_226_I8_carry_5_port, S => 
                           position1_N2306);
   position1_sub_226_I8_U2_5 : ADD32 port map( A => n933, B => n42, CI => 
                           position1_sub_226_I8_carry_5_port, CO => 
                           position1_sub_226_I8_carry_6_port, S => 
                           position1_N2307);
   position1_sub_226_I8_U2_6 : ADD32 port map( A => n932, B => n250, CI => 
                           position1_sub_226_I8_carry_6_port, CO => 
                           position1_sub_226_I8_carry_7_port, S => 
                           position1_N2308);
   position1_sub_226_I8_U2_7 : ADD32 port map( A => n930, B => n46, CI => 
                           position1_sub_226_I8_carry_7_port, CO => 
                           position1_sub_226_I8_carry_8_port, S => 
                           position1_N2309);
   position1_sub_226_I8_U2_8 : ADD32 port map( A => n929, B => n254, CI => 
                           position1_sub_226_I8_carry_8_port, CO => 
                           position1_sub_226_I8_carry_9_port, S => 
                           position1_N2310);
   position1_sub_226_I8_U2_9 : ADD32 port map( A => n927, B => n41, CI => 
                           position1_sub_226_I8_carry_9_port, CO => 
                           position1_sub_226_I8_carry_10_port, S => 
                           position1_N2311);
   position1_sub_226_I8_U2_10 : ADD32 port map( A => n926, B => n286, CI => 
                           position1_sub_226_I8_carry_10_port, CO => 
                           position1_sub_226_I8_carry_11_port, S => 
                           position1_N2312);
   position1_sub_226_I8_U2_11 : ADD32 port map( A => n925, B => n47, CI => 
                           position1_sub_226_I8_carry_11_port, CO => 
                           position1_sub_226_I8_carry_12_port, S => 
                           position1_N2313);
   position1_sub_226_I8_U2_12 : ADD32 port map( A => n923, B => n290, CI => 
                           position1_sub_226_I8_carry_12_port, CO => 
                           position1_sub_226_I8_carry_13_port, S => 
                           position1_N2314);
   position1_sub_226_I8_U2_13 : ADD32 port map( A => n921, B => n44, CI => 
                           position1_sub_226_I8_carry_13_port, CO => 
                           position1_sub_226_I8_carry_14_port, S => 
                           position1_N2315);
   position1_sub_226_I8_U2_14 : ADD32 port map( A => n920, B => n294, CI => 
                           position1_sub_226_I8_carry_14_port, CO => 
                           position1_sub_226_I8_carry_15_port, S => 
                           position1_N2316);
   position1_sub_226_I8_U2_15 : ADD32 port map( A => n918, B => n43, CI => 
                           position1_sub_226_I8_carry_15_port, CO => 
                           position1_sub_226_I8_carry_16_port, S => 
                           position1_N2317);
   position1_sub_226_I8_U2_16 : ADD32 port map( A => n917, B => n298, CI => 
                           position1_sub_226_I8_carry_16_port, CO => 
                           position1_sub_226_I8_carry_17_port, S => 
                           position1_N2318);
   position1_sub_226_I8_U2_17 : ADD32 port map( A => n916, B => n45, CI => 
                           position1_sub_226_I8_carry_17_port, CO => 
                           position1_sub_226_I8_carry_18_port, S => 
                           position1_N2319);
   position1_sub_226_I8_U2_18 : ADD32 port map( A => n915, B => n592, CI => 
                           position1_sub_226_I8_carry_18_port, CO => 
                           position1_sub_226_I8_carry_19_port, S => 
                           position1_N2320);
   position1_dp_cluster_0_add_196_aco_U1_1 : ADD32 port map( A => 
                           position1_x_sum_1_port, B => n837, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_1_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_2_port, 
                           S => position1_N1178_port);
   position1_dp_cluster_0_add_196_aco_U1_2 : ADD32 port map( A => 
                           position1_x_sum_2_port, B => n857, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_2_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_3_port, 
                           S => position1_N1179_port);
   position1_dp_cluster_0_add_196_aco_U1_3 : ADD32 port map( A => 
                           position1_x_sum_3_port, B => n859, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_3_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_4_port, 
                           S => position1_N1180_port);
   position1_dp_cluster_0_add_196_aco_U1_4 : ADD32 port map( A => 
                           position1_x_sum_4_port, B => n861, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_4_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_5_port, 
                           S => position1_N1181_port);
   position1_dp_cluster_0_add_196_aco_U1_5 : ADD32 port map( A => 
                           position1_x_sum_5_port, B => n863, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_5_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_6_port, 
                           S => position1_N1182_port);
   position1_dp_cluster_0_add_196_aco_U1_6 : ADD32 port map( A => 
                           position1_x_sum_6_port, B => n865, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_6_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_7_port, 
                           S => position1_N1183_port);
   position1_dp_cluster_0_add_196_aco_U1_7 : ADD32 port map( A => 
                           position1_x_sum_7_port, B => n868, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_7_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_8_port, 
                           S => position1_N1184_port);
   position1_dp_cluster_0_add_196_aco_U1_8 : ADD32 port map( A => 
                           position1_x_sum_8_port, B => n870, CI => 
                           position1_dp_cluster_0_add_196_aco_carry_8_port, CO 
                           => position1_dp_cluster_0_add_196_aco_carry_9_port, 
                           S => position1_N1185_port);
   position1_dp_cluster_1_add_197_aco_U1_1 : ADD32 port map( A => 
                           position1_y_sum_1_port, B => n810, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_1_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_2_port, 
                           S => position1_N1203_port);
   position1_dp_cluster_1_add_197_aco_U1_2 : ADD32 port map( A => 
                           position1_y_sum_2_port, B => n806, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_2_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_3_port, 
                           S => position1_N1204_port);
   position1_dp_cluster_1_add_197_aco_U1_3 : ADD32 port map( A => 
                           position1_y_sum_3_port, B => n802, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_3_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_4_port, 
                           S => position1_N1205_port);
   position1_dp_cluster_1_add_197_aco_U1_4 : ADD32 port map( A => 
                           position1_y_sum_4_port, B => n798, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_4_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_5_port, 
                           S => position1_N1206_port);
   position1_dp_cluster_1_add_197_aco_U1_5 : ADD32 port map( A => 
                           position1_y_sum_5_port, B => n794, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_5_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_6_port, 
                           S => position1_N1207_port);
   position1_dp_cluster_1_add_197_aco_U1_6 : ADD32 port map( A => 
                           position1_y_sum_6_port, B => n790, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_6_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_7_port, 
                           S => position1_N1208_port);
   position1_dp_cluster_1_add_197_aco_U1_7 : ADD32 port map( A => 
                           position1_y_sum_7_port, B => n786, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_7_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_8_port, 
                           S => position1_N1209_port);
   position1_dp_cluster_1_add_197_aco_U1_8 : ADD32 port map( A => 
                           position1_y_sum_8_port, B => n780, CI => 
                           position1_dp_cluster_1_add_197_aco_carry_8_port, CO 
                           => position1_dp_cluster_1_add_197_aco_carry_9_port, 
                           S => position1_N1210_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_2 : ADD32 port map( A => 
                           position1_N357_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_2_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_3_port, S 
                           => position1_N981_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_3 : ADD32 port map( A => 
                           position1_N358_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_3_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_4_port, S 
                           => position1_N982_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_4 : ADD32 port map( A => 
                           position1_N359, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_4_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_5_port, S 
                           => position1_N983_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_5 : ADD32 port map( A => 
                           position1_N360_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_5_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_6_port, S 
                           => position1_N984_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_6 : ADD32 port map( A => 
                           position1_N361, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_6_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_7_port, S 
                           => position1_N985_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_7 : ADD32 port map( A => 
                           position1_N362_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_7_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_8_port, S 
                           => position1_N986_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_8 : ADD32 port map( A => 
                           position1_N363_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, 
                           CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_8_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_9_port, S 
                           => position1_N987_port);
   position1_dp_cluster_2_add_0_root_add_189_3_U1_9 : ADD32 port map( A => 
                           position1_N364_port, B => 
                           position1_dp_cluster_6_N389, CI => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_9_port, 
                           CO => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_10_port, S 
                           => position1_N988_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_2 : ADD32 port map( A => 
                           position1_N282, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_2_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_2_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_3_port, S 
                           => position1_N906_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_3 : ADD32 port map( A => 
                           position1_N283_port, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_3_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_3_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_4_port, S 
                           => position1_N907_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_4 : ADD32 port map( A => 
                           position1_N284, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_4_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_4_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_5_port, S 
                           => position1_N908_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_5 : ADD32 port map( A => 
                           position1_N285, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_5_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_5_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_6_port, S 
                           => position1_N909_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_6 : ADD32 port map( A => 
                           position1_N286, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_6_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_6_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_7_port, S 
                           => position1_N910_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_7 : ADD32 port map( A => 
                           position1_N287, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_7_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_7_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_8_port, S 
                           => position1_N911_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_8 : ADD32 port map( A => 
                           position1_N288, B => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_8_port, 
                           CI => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_8_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_9_port, S 
                           => position1_N912_port);
   position1_dp_cluster_3_add_0_root_add_188_3_U1_9 : ADD32 port map( A => 
                           position1_N289, B => position1_dp_cluster_7_N314, CI
                           => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_9_port, 
                           CO => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_10_port, S 
                           => position1_N913_port);
   position1_dp_cluster_4_add_178_aco_U1_1 : ADD32 port map( A => 
                           position1_x_sum_1_port, B => n836, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_1_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_2_port, 
                           S => position1_N608);
   position1_dp_cluster_4_add_178_aco_U1_2 : ADD32 port map( A => 
                           position1_x_sum_2_port, B => n856, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_2_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_3_port, 
                           S => position1_N609);
   position1_dp_cluster_4_add_178_aco_U1_3 : ADD32 port map( A => 
                           position1_x_sum_3_port, B => n858, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_3_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_4_port, 
                           S => position1_N610);
   position1_dp_cluster_4_add_178_aco_U1_4 : ADD32 port map( A => 
                           position1_x_sum_4_port, B => n860, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_4_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_5_port, 
                           S => position1_N611);
   position1_dp_cluster_4_add_178_aco_U1_5 : ADD32 port map( A => 
                           position1_x_sum_5_port, B => n862, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_5_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_6_port, 
                           S => position1_N612);
   position1_dp_cluster_4_add_178_aco_U1_6 : ADD32 port map( A => 
                           position1_x_sum_6_port, B => n864, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_6_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_7_port, 
                           S => position1_N613);
   position1_dp_cluster_4_add_178_aco_U1_7 : ADD32 port map( A => 
                           position1_x_sum_7_port, B => n867, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_7_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_8_port, 
                           S => position1_N614);
   position1_dp_cluster_4_add_178_aco_U1_8 : ADD32 port map( A => 
                           position1_x_sum_8_port, B => n869, CI => 
                           position1_dp_cluster_4_add_178_aco_carry_8_port, CO 
                           => position1_dp_cluster_4_add_178_aco_carry_9_port, 
                           S => position1_N615);
   position1_dp_cluster_5_add_179_aco_U1_1 : ADD32 port map( A => 
                           position1_y_sum_1_port, B => n809, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_1_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_2_port, 
                           S => position1_N633);
   position1_dp_cluster_5_add_179_aco_U1_2 : ADD32 port map( A => 
                           position1_y_sum_2_port, B => n805, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_2_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_3_port, 
                           S => position1_N634);
   position1_dp_cluster_5_add_179_aco_U1_3 : ADD32 port map( A => 
                           position1_y_sum_3_port, B => n801, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_3_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_4_port, 
                           S => position1_N635);
   position1_dp_cluster_5_add_179_aco_U1_4 : ADD32 port map( A => 
                           position1_y_sum_4_port, B => n797, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_4_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_5_port, 
                           S => position1_N636);
   position1_dp_cluster_5_add_179_aco_U1_5 : ADD32 port map( A => 
                           position1_y_sum_5_port, B => n793, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_5_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_6_port, 
                           S => position1_N637);
   position1_dp_cluster_5_add_179_aco_U1_6 : ADD32 port map( A => 
                           position1_y_sum_6_port, B => n789, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_6_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_7_port, 
                           S => position1_N638);
   position1_dp_cluster_5_add_179_aco_U1_7 : ADD32 port map( A => 
                           position1_y_sum_7_port, B => n785, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_7_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_8_port, 
                           S => position1_N639);
   position1_dp_cluster_5_add_179_aco_U1_8 : ADD32 port map( A => 
                           position1_y_sum_8_port, B => n779, CI => 
                           position1_dp_cluster_5_add_179_aco_carry_8_port, CO 
                           => position1_dp_cluster_5_add_179_aco_carry_9_port, 
                           S => position1_N640);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_2 : ADD32 port map( A => 
                           position1_N357_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_2_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_3_port, S 
                           => position1_N407);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_3 : ADD32 port map( A => 
                           position1_N358_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_3_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_4_port, S 
                           => position1_N408);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_4 : ADD32 port map( A => 
                           position1_N359, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_4_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_5_port, S 
                           => position1_N409);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_5 : ADD32 port map( A => 
                           position1_N360_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_5_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_6_port, S 
                           => position1_N410);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_6 : ADD32 port map( A => 
                           position1_N361, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_6_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_7_port, S 
                           => position1_N411);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_7 : ADD32 port map( A => 
                           position1_N362_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_7_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_8_port, S 
                           => position1_N412);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_8 : ADD32 port map( A => 
                           position1_N363_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, 
                           CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_8_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_9_port, S 
                           => position1_N413);
   position1_dp_cluster_6_add_0_root_add_171_3_U1_9 : ADD32 port map( A => 
                           position1_N364_port, B => 
                           position1_dp_cluster_6_N389, CI => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_9_port, 
                           CO => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_10_port, S 
                           => position1_N414);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_2 : ADD32 port map( A => 
                           position1_N282, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_2_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_2_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_3_port, S 
                           => position1_N332);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_3 : ADD32 port map( A => 
                           position1_N283_port, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_3_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_3_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_4_port, S 
                           => position1_N333);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_4 : ADD32 port map( A => 
                           position1_N284, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_4_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_4_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_5_port, S 
                           => position1_N334);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_5 : ADD32 port map( A => 
                           position1_N285, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_5_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_5_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_6_port, S 
                           => position1_N335);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_6 : ADD32 port map( A => 
                           position1_N286, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_6_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_6_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_7_port, S 
                           => position1_N336);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_7 : ADD32 port map( A => 
                           position1_N287, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_7_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_7_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_8_port, S 
                           => position1_N337);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_8 : ADD32 port map( A => 
                           position1_N288, B => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_8_port, 
                           CI => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_8_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_9_port, S 
                           => position1_N338);
   position1_dp_cluster_7_add_0_root_add_170_3_U1_9 : ADD32 port map( A => 
                           position1_N289, B => position1_dp_cluster_7_N314, CI
                           => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_9_port, 
                           CO => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_10_port, S 
                           => position1_N339);
   gensync1_add_39_U1_1_1 : ADD22 port map( A => gensync1_N182, B => 
                           gensync1_N74, CO => gensync1_add_39_carry_2_port, S 
                           => gensync1_N13);
   gensync1_add_39_U1_1_2 : ADD22 port map( A => gensync1_N181, B => 
                           gensync1_add_39_carry_2_port, CO => 
                           gensync1_add_39_carry_3_port, S => gensync1_N14);
   gensync1_add_39_U1_1_3 : ADD22 port map( A => gensync1_N180, B => 
                           gensync1_add_39_carry_3_port, CO => 
                           gensync1_add_39_carry_4_port, S => gensync1_N15);
   gensync1_add_39_U1_1_4 : ADD22 port map( A => gensync1_N179, B => 
                           gensync1_add_39_carry_4_port, CO => 
                           gensync1_add_39_carry_5_port, S => gensync1_N16);
   gensync1_add_39_U1_1_5 : ADD22 port map( A => gensync1_N178, B => 
                           gensync1_add_39_carry_5_port, CO => 
                           gensync1_add_39_carry_6_port, S => gensync1_N17);
   gensync1_add_39_U1_1_6 : ADD22 port map( A => gensync1_N177, B => 
                           gensync1_add_39_carry_6_port, CO => 
                           gensync1_add_39_carry_7_port, S => gensync1_N18);
   gensync1_add_39_U1_1_7 : ADD22 port map( A => gensync1_N176, B => 
                           gensync1_add_39_carry_7_port, CO => 
                           gensync1_add_39_carry_8_port, S => gensync1_N19);
   gensync1_add_39_U1_1_8 : ADD22 port map( A => n477, B => 
                           gensync1_add_39_carry_8_port, CO => 
                           gensync1_add_39_carry_9_port, S => gensync1_N20);
   gensync1_add_45_U1_1_1 : ADD22 port map( A => gensync1_N172, B => 
                           gensync1_N173, CO => gensync1_add_45_carry_2_port, S
                           => gensync1_N47);
   gensync1_add_45_U1_1_2 : ADD22 port map( A => gensync1_N171, B => 
                           gensync1_add_45_carry_2_port, CO => 
                           gensync1_add_45_carry_3_port, S => gensync1_N48);
   gensync1_add_45_U1_1_3 : ADD22 port map( A => gensync1_N170, B => 
                           gensync1_add_45_carry_3_port, CO => 
                           gensync1_add_45_carry_4_port, S => gensync1_N49);
   gensync1_add_45_U1_1_4 : ADD22 port map( A => gensync1_N169, B => 
                           gensync1_add_45_carry_4_port, CO => 
                           gensync1_add_45_carry_5_port, S => gensync1_N50);
   gensync1_add_45_U1_1_5 : ADD22 port map( A => gensync1_N168, B => 
                           gensync1_add_45_carry_5_port, CO => 
                           gensync1_add_45_carry_6_port, S => gensync1_N51);
   gensync1_add_45_U1_1_6 : ADD22 port map( A => gensync1_N167, B => 
                           gensync1_add_45_carry_6_port, CO => 
                           gensync1_add_45_carry_7_port, S => gensync1_N52);
   gensync1_add_45_U1_1_7 : ADD22 port map( A => gensync1_N166, B => 
                           gensync1_add_45_carry_7_port, CO => 
                           gensync1_add_45_carry_8_port, S => gensync1_N53);
   gensync1_add_45_U1_1_8 : ADD22 port map( A => gensync1_N165, B => 
                           gensync1_add_45_carry_8_port, CO => 
                           gensync1_add_45_carry_9_port, S => gensync1_N54);
   gensync1_VSYNC_reg : DF3 port map( D => n817, C => CLK_top, Q => VSYNC_top, 
                           QN => n_1000);
   gensync1_HSYNC_reg : DF3 port map( D => n874, C => CLK_top, Q => HSYNC_top, 
                           QN => n_1001);
   gensync1_comptX_reg_1_inst : DF3 port map( D => gensync1_N23, C => CLK_top, 
                           Q => gensync1_N182, QN => n10);
   gensync1_comptX_reg_2_inst : DF3 port map( D => gensync1_N24, C => CLK_top, 
                           Q => gensync1_N181, QN => n4);
   gensync1_comptX_reg_3_inst : DF3 port map( D => gensync1_N25, C => CLK_top, 
                           Q => gensync1_N180, QN => n12);
   gensync1_comptX_reg_4_inst : DF3 port map( D => gensync1_N26, C => CLK_top, 
                           Q => gensync1_N179, QN => n7);
   gensync1_comptX_reg_5_inst : DF3 port map( D => gensync1_N27, C => CLK_top, 
                           Q => gensync1_N178, QN => n14);
   gensync1_comptX_reg_6_inst : DF3 port map( D => gensync1_N28, C => CLK_top, 
                           Q => gensync1_N177, QN => n6);
   gensync1_comptX_reg_7_inst : DF3 port map( D => gensync1_N29, C => CLK_top, 
                           Q => gensync1_N176, QN => n15);
   gensync1_comptX_reg_8_inst : DF3 port map( D => gensync1_N30, C => CLK_top, 
                           Q => gensync1_N175, QN => n_1002);
   gensync1_comptX_reg_9_inst : DF3 port map( D => gensync1_N31, C => CLK_top, 
                           Q => gensync1_N174, QN => n_1003);
   gensync1_comptX_reg_0_inst : DF3 port map( D => gensync1_N22, C => CLK_top, 
                           Q => gensync1_N74, QN => n1);
   image_process1_state_reg : DF3 port map( D => reset_top, C => CLK_top, Q => 
                           image_process1_state, QN => image_process1_n27);
   image_process1_bi_reg_0_inst : DF3 port map( D => n751, C => CLK_top, Q => 
                           image_process1_bi_0_port, QN => n_1004);
   image_process1_bi_reg_1_inst : DF3 port map( D => n750, C => CLK_top, Q => 
                           image_process1_bi_1_port, QN => n_1005);
   image_process1_bi_reg_2_inst : DF3 port map( D => n749, C => CLK_top, Q => 
                           n_1006, QN => image_process1_n25);
   image_process1_bi_reg_3_inst : DF3 port map( D => n748, C => CLK_top, Q => 
                           image_process1_bi_3_port, QN => n_1007);
   image_process1_bi_reg_4_inst : DF3 port map( D => n747, C => CLK_top, Q => 
                           image_process1_bi_4_port, QN => n_1008);
   image_process1_bi_reg_5_inst : DF3 port map( D => n746, C => CLK_top, Q => 
                           image_process1_bi_5_port, QN => n_1009);
   image_process1_bi_reg_6_inst : DF3 port map( D => n745, C => CLK_top, Q => 
                           image_process1_bi_6_port, QN => n_1010);
   image_process1_bi_reg_7_inst : DF3 port map( D => n744, C => CLK_top, Q => 
                           image_process1_bi_7_port, QN => n_1011);
   image_process1_gi_reg_0_inst : DF3 port map( D => n759, C => CLK_top, Q => 
                           image_process1_gi_0_port, QN => n_1012);
   image_process1_gi_reg_1_inst : DF3 port map( D => n758, C => CLK_top, Q => 
                           image_process1_gi_1_port, QN => n_1013);
   image_process1_gi_reg_2_inst : DF3 port map( D => n757, C => CLK_top, Q => 
                           image_process1_gi_2_port, QN => n_1014);
   image_process1_gi_reg_3_inst : DF3 port map( D => n756, C => CLK_top, Q => 
                           image_process1_gi_3_port, QN => n_1015);
   image_process1_gi_reg_4_inst : DF3 port map( D => n755, C => CLK_top, Q => 
                           image_process1_gi_4_port, QN => n5);
   image_process1_gi_reg_5_inst : DF3 port map( D => n754, C => CLK_top, Q => 
                           image_process1_gi_5_port, QN => n33);
   image_process1_gi_reg_6_inst : DF3 port map( D => n753, C => CLK_top, Q => 
                           image_process1_gi_6_port, QN => n_1016);
   image_process1_gi_reg_7_inst : DF3 port map( D => n752, C => CLK_top, Q => 
                           image_process1_gi_7_port, QN => n_1017);
   image_process1_ri_reg_0_inst : DF3 port map( D => n767, C => CLK_top, Q => 
                           image_process1_ri_0_port, QN => n_1018);
   image_process1_ri_reg_1_inst : DF3 port map( D => n766, C => CLK_top, Q => 
                           image_process1_ri_1_port, QN => n_1019);
   image_process1_ri_reg_2_inst : DF3 port map( D => n765, C => CLK_top, Q => 
                           n_1020, QN => image_process1_n13);
   image_process1_ri_reg_3_inst : DF3 port map( D => n764, C => CLK_top, Q => 
                           image_process1_ri_3_port, QN => n_1021);
   image_process1_ri_reg_4_inst : DF3 port map( D => n763, C => CLK_top, Q => 
                           image_process1_ri_4_port, QN => n_1022);
   image_process1_ri_reg_5_inst : DF3 port map( D => n762, C => CLK_top, Q => 
                           image_process1_ri_5_port, QN => n_1023);
   image_process1_ri_reg_6_inst : DF3 port map( D => n761, C => CLK_top, Q => 
                           image_process1_ri_6_port, QN => n_1024);
   image_process1_ri_reg_7_inst : DF3 port map( D => n760, C => CLK_top, Q => 
                           image_process1_ri_7_port, QN => n_1025);
   position1_b_bout_reg_3_inst : DF3 port map( D => position1_N100, C => 
                           CLK_top, Q => bout_top(3), QN => n_1026);
   position1_b_bout_reg_4_inst : DF3 port map( D => position1_N101, C => 
                           CLK_top, Q => bout_top(4), QN => n_1027);
   position1_b_bout_reg_5_inst : DF3 port map( D => position1_N102, C => 
                           CLK_top, Q => bout_top(5), QN => n_1028);
   position1_b_bout_reg_6_inst : DF3 port map( D => position1_N103, C => 
                           CLK_top, Q => bout_top(6), QN => n_1029);
   position1_b_bout_reg_7_inst : DF3 port map( D => position1_N104, C => 
                           CLK_top, Q => bout_top(7), QN => n_1030);
   position1_r_bout_reg_0_inst : DF3 port map( D => position1_N81, C => CLK_top
                           , Q => rout_top(0), QN => n_1031);
   position1_r_bout_reg_1_inst : DF3 port map( D => position1_N82, C => CLK_top
                           , Q => rout_top(1), QN => n_1032);
   position1_r_bout_reg_2_inst : DF3 port map( D => position1_N83, C => CLK_top
                           , Q => rout_top(2), QN => n_1033);
   position1_r_bout_reg_3_inst : DF3 port map( D => position1_N84, C => CLK_top
                           , Q => rout_top(3), QN => n_1034);
   position1_r_bout_reg_4_inst : DF3 port map( D => position1_N85, C => CLK_top
                           , Q => rout_top(4), QN => n_1035);
   position1_r_bout_reg_5_inst : DF3 port map( D => position1_N86, C => CLK_top
                           , Q => rout_top(5), QN => n_1036);
   position1_r_bout_reg_6_inst : DF3 port map( D => position1_N87, C => CLK_top
                           , Q => rout_top(6), QN => n_1037);
   position1_r_bout_reg_7_inst : DF3 port map( D => position1_N88, C => CLK_top
                           , Q => rout_top(7), QN => n_1038);
   position1_b_bout_reg_0_inst : DF3 port map( D => position1_N97, C => CLK_top
                           , Q => bout_top(0), QN => n_1039);
   position1_b_bout_reg_1_inst : DF3 port map( D => position1_N98, C => CLK_top
                           , Q => bout_top(1), QN => n_1040);
   position1_b_bout_reg_2_inst : DF3 port map( D => position1_N99, C => CLK_top
                           , Q => bout_top(2), QN => n_1041);
   position1_g_bout_reg_1_inst : DF3 port map( D => n715, C => CLK_top, Q => 
                           gout_top(1), QN => n_1042);
   position1_g_bout_reg_3_inst : DF3 port map( D => n716, C => CLK_top, Q => 
                           gout_top(3), QN => n_1043);
   position1_g_bout_reg_7_inst : DF3 port map( D => n717, C => CLK_top, Q => 
                           gout_top(7), QN => n_1044);
   position1_g_bout_reg_0_inst : DF3 port map( D => position1_N89, C => CLK_top
                           , Q => gout_top(0), QN => n_1045);
   position1_g_bout_reg_2_inst : DF3 port map( D => position1_N91, C => CLK_top
                           , Q => gout_top(2), QN => n_1046);
   position1_g_bout_reg_4_inst : DF3 port map( D => position1_N93, C => CLK_top
                           , Q => gout_top(4), QN => n_1047);
   position1_g_bout_reg_5_inst : DF3 port map( D => position1_N94, C => CLK_top
                           , Q => gout_top(5), QN => n_1048);
   position1_g_bout_reg_6_inst : DF3 port map( D => position1_N95, C => CLK_top
                           , Q => gout_top(6), QN => n_1049);
   position1_y_bar_reg_0_inst : DF3 port map( D => n685, C => CLK_top, Q => 
                           Y_barycentre_top_0_port, QN => n_1050);
   position1_quot_y_reg_0_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2363, GN => n1360, Q => 
                           position1_quot_y_0_port);
   position1_y_bar_reg_1_inst : DF3 port map( D => n686, C => CLK_top, Q => 
                           Y_barycentre_top_1_port, QN => n23);
   position1_quot_y_reg_1_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2364, GN => n1360, Q => 
                           position1_quot_y_1_port);
   position1_y_bar_reg_2_inst : DF3 port map( D => n687, C => CLK_top, Q => 
                           Y_barycentre_top_2_port, QN => n21);
   position1_quot_y_reg_2_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2365, GN => n1360, Q => 
                           position1_quot_y_2_port);
   position1_y_bar_reg_3_inst : DF3 port map( D => n688, C => CLK_top, Q => 
                           Y_barycentre_top_3_port, QN => n24);
   position1_quot_y_reg_3_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2366, GN => n1360, Q => 
                           position1_quot_y_3_port);
   position1_y_bar_reg_4_inst : DF3 port map( D => n689, C => CLK_top, Q => 
                           Y_barycentre_top_4_port, QN => n26);
   position1_quot_y_reg_4_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2367, GN => n1360, Q => 
                           position1_quot_y_4_port);
   position1_y_bar_reg_5_inst : DF3 port map( D => n690, C => CLK_top, Q => 
                           Y_barycentre_top_5_port, QN => n28);
   position1_quot_y_reg_5_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2368, GN => n1360, Q => 
                           position1_quot_y_5_port);
   position1_y_bar_reg_6_inst : DF3 port map( D => n691, C => CLK_top, Q => 
                           Y_barycentre_top_6_port, QN => n31);
   position1_quot_y_reg_6_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2369, GN => n1360, Q => 
                           position1_quot_y_6_port);
   position1_y_bar_reg_7_inst : DF3 port map( D => n692, C => CLK_top, Q => 
                           Y_barycentre_top_7_port, QN => n32);
   position1_quot_y_reg_7_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2370, GN => n1360, Q => 
                           position1_quot_y_7_port);
   position1_y_bar_reg_8_inst : DF3 port map( D => n693, C => CLK_top, Q => 
                           Y_barycentre_top_8_port, QN => n30);
   position1_quot_y_reg_8_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2371, GN => n1360, Q => 
                           position1_quot_y_8_port);
   position1_x_bar_reg_0_inst : DF3 port map( D => n676, C => CLK_top, Q => 
                           X_barycentre_top_0_port, QN => n_1051);
   position1_quot_x_reg_0_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2354, GN => n1360, Q => 
                           position1_quot_x_0_port);
   position1_x_bar_reg_1_inst : DF3 port map( D => n677, C => CLK_top, Q => 
                           X_barycentre_top_1_port, QN => n17);
   position1_quot_x_reg_1_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2355, GN => n1360, Q => 
                           position1_quot_x_1_port);
   position1_x_bar_reg_2_inst : DF3 port map( D => n678, C => CLK_top, Q => 
                           X_barycentre_top_2_port, QN => n16);
   position1_quot_x_reg_2_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2356, GN => n1360, Q => 
                           position1_quot_x_2_port);
   position1_x_bar_reg_3_inst : DF3 port map( D => n679, C => CLK_top, Q => 
                           X_barycentre_top_3_port, QN => n19);
   position1_quot_x_reg_3_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2357, GN => n1360, Q => 
                           position1_quot_x_3_port);
   position1_x_bar_reg_4_inst : DF3 port map( D => n680, C => CLK_top, Q => 
                           X_barycentre_top_4_port, QN => n20);
   position1_quot_x_reg_4_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2358, GN => n1360, Q => 
                           position1_quot_x_4_port);
   position1_x_bar_reg_5_inst : DF3 port map( D => n681, C => CLK_top, Q => 
                           X_barycentre_top_5_port, QN => n22);
   position1_quot_x_reg_5_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2359, GN => n1360, Q => 
                           position1_quot_x_5_port);
   position1_x_bar_reg_6_inst : DF3 port map( D => n682, C => CLK_top, Q => 
                           X_barycentre_top_6_port, QN => n25);
   position1_quot_x_reg_6_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2360, GN => n1360, Q => 
                           position1_quot_x_6_port);
   position1_x_bar_reg_7_inst : DF3 port map( D => n683, C => CLK_top, Q => 
                           X_barycentre_top_7_port, QN => n27);
   position1_quot_x_reg_7_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2361, GN => n1360, Q => 
                           position1_quot_x_7_port);
   position1_x_bar_reg_8_inst : DF3 port map( D => n684, C => CLK_top, Q => 
                           X_barycentre_top_8_port, QN => n29);
   position1_quot_x_reg_8_inst : DLPQ3 port map( SN => position1_n283, D => 
                           position1_N2362, GN => n1360, Q => 
                           position1_quot_x_8_port);
   position1_count_reg_15_inst : DF3 port map( D => n672, C => CLK_top, Q => 
                           position1_N2446, QN => n68);
   position1_count_reg_14_inst : DF3 port map( D => n671, C => CLK_top, Q => 
                           position1_N2447, QN => n43);
   position1_count_reg_13_inst : DF3 port map( D => n670, C => CLK_top, Q => 
                           position1_N2448, QN => n40);
   position1_count_reg_12_inst : DF3 port map( D => n669, C => CLK_top, Q => 
                           position1_N2449, QN => n44);
   position1_count_reg_11_inst : DF3 port map( D => n668, C => CLK_top, Q => 
                           position1_N2450, QN => n39);
   position1_count_reg_10_inst : DF3 port map( D => n667, C => CLK_top, Q => 
                           position1_N2451, QN => n47);
   position1_count_reg_9_inst : DF3 port map( D => n666, C => CLK_top, Q => 
                           position1_N2452, QN => n36);
   position1_count_reg_8_inst : DF3 port map( D => n665, C => CLK_top, Q => 
                           position1_N2453, QN => n41);
   position1_count_reg_7_inst : DF3 port map( D => n664, C => CLK_top, Q => 
                           position1_N2454, QN => n101);
   position1_count_reg_6_inst : DF3 port map( D => n663, C => CLK_top, Q => 
                           position1_N2455, QN => n46);
   position1_count_reg_5_inst : DF3 port map( D => n662, C => CLK_top, Q => 
                           position1_N2456, QN => n48);
   position1_count_reg_4_inst : DF3 port map( D => n661, C => CLK_top, Q => 
                           position1_N2457, QN => n42);
   position1_count_reg_3_inst : DF3 port map( D => n660, C => CLK_top, Q => 
                           position1_N2458, QN => n38);
   position1_count_reg_2_inst : DF3 port map( D => n659, C => CLK_top, Q => 
                           position1_N2459, QN => n67);
   position1_count_reg_1_inst : DF3 port map( D => n658, C => CLK_top, Q => 
                           position1_N2460, QN => n37);
   position1_count_reg_16_inst : DF3 port map( D => n673, C => CLK_top, Q => 
                           position1_N2445, QN => n45);
   position1_count_reg_17_inst : DF3 port map( D => n674, C => CLK_top, Q => n2
                           , QN => n102);
   position1_count_reg_0_inst : DF3 port map( D => n657, C => CLK_top, Q => 
                           position1_N560, QN => n35);
   position1_x_sum_reg_22_inst : DF3 port map( D => position1_n1613, C => 
                           CLK_top, Q => position1_x_sum_22_port, QN => n77);
   position1_x_sum_reg_21_inst : DF3 port map( D => position1_n1614, C => 
                           CLK_top, Q => position1_x_sum_21_port, QN => n61);
   position1_x_sum_reg_20_inst : DF3 port map( D => position1_n1615, C => 
                           CLK_top, Q => position1_x_sum_20_port, QN => n78);
   position1_x_sum_reg_19_inst : DF3 port map( D => position1_n1616, C => 
                           CLK_top, Q => position1_x_sum_19_port, QN => n62);
   position1_x_sum_reg_18_inst : DF3 port map( D => position1_n1617, C => 
                           CLK_top, Q => position1_x_sum_18_port, QN => n79);
   position1_x_sum_reg_17_inst : DF3 port map( D => position1_n1618, C => 
                           CLK_top, Q => position1_x_sum_17_port, QN => n63);
   position1_x_sum_reg_16_inst : DF3 port map( D => position1_n1619, C => 
                           CLK_top, Q => position1_x_sum_16_port, QN => n80);
   position1_x_sum_reg_15_inst : DF3 port map( D => position1_n1620, C => 
                           CLK_top, Q => position1_x_sum_15_port, QN => n64);
   position1_x_sum_reg_14_inst : DF3 port map( D => position1_n1621, C => 
                           CLK_top, Q => position1_x_sum_14_port, QN => n81);
   position1_x_sum_reg_13_inst : DF3 port map( D => position1_n1622, C => 
                           CLK_top, Q => position1_x_sum_13_port, QN => n65);
   position1_x_sum_reg_12_inst : DF3 port map( D => position1_n1623, C => 
                           CLK_top, Q => position1_x_sum_12_port, QN => n82);
   position1_x_sum_reg_11_inst : DF3 port map( D => position1_n1624, C => 
                           CLK_top, Q => position1_x_sum_11_port, QN => n66);
   position1_x_sum_reg_10_inst : DF3 port map( D => position1_n1625, C => 
                           CLK_top, Q => position1_x_sum_10_port, QN => n70);
   position1_x_sum_reg_9_inst : DF3 port map( D => position1_n1626, C => 
                           CLK_top, Q => position1_x_sum_9_port, QN => n52);
   position1_x_sum_reg_8_inst : DF3 port map( D => position1_n1627, C => 
                           CLK_top, Q => position1_x_sum_8_port, QN => n50);
   position1_x_sum_reg_7_inst : DF3 port map( D => position1_n1628, C => 
                           CLK_top, Q => position1_x_sum_7_port, QN => n95);
   position1_x_sum_reg_6_inst : DF3 port map( D => position1_n1629, C => 
                           CLK_top, Q => position1_x_sum_6_port, QN => n88);
   position1_x_sum_reg_5_inst : DF3 port map( D => position1_n1630, C => 
                           CLK_top, Q => position1_x_sum_5_port, QN => n89);
   position1_x_sum_reg_4_inst : DF3 port map( D => position1_n1631, C => 
                           CLK_top, Q => position1_x_sum_4_port, QN => n90);
   position1_x_sum_reg_3_inst : DF3 port map( D => position1_n1632, C => 
                           CLK_top, Q => position1_x_sum_3_port, QN => n96);
   position1_x_sum_reg_2_inst : DF3 port map( D => position1_n1633, C => 
                           CLK_top, Q => position1_x_sum_2_port, QN => n91);
   position1_x_sum_reg_1_inst : DF3 port map( D => position1_n1634, C => 
                           CLK_top, Q => position1_x_sum_1_port, QN => n92);
   position1_x_sum_reg_23_inst : DF3 port map( D => position1_n1612, C => 
                           CLK_top, Q => position1_x_sum_23_port, QN => n60);
   position1_x_sum_reg_24_inst : DF3 port map( D => position1_n1611, C => 
                           CLK_top, Q => position1_x_sum_24_port, QN => n100);
   position1_x_sum_reg_0_inst : DF3 port map( D => position1_n1635, C => 
                           CLK_top, Q => position1_N1521_port, QN => n98);
   position1_y_sum_reg_22_inst : DF3 port map( D => position1_n1588, C => 
                           CLK_top, Q => position1_y_sum_22_port, QN => n71);
   position1_y_sum_reg_21_inst : DF3 port map( D => position1_n1589, C => 
                           CLK_top, Q => position1_y_sum_21_port, QN => n54);
   position1_y_sum_reg_20_inst : DF3 port map( D => position1_n1590, C => 
                           CLK_top, Q => position1_y_sum_20_port, QN => n72);
   position1_y_sum_reg_19_inst : DF3 port map( D => position1_n1591, C => 
                           CLK_top, Q => position1_y_sum_19_port, QN => n55);
   position1_y_sum_reg_18_inst : DF3 port map( D => position1_n1592, C => 
                           CLK_top, Q => position1_y_sum_18_port, QN => n73);
   position1_y_sum_reg_17_inst : DF3 port map( D => position1_n1593, C => 
                           CLK_top, Q => position1_y_sum_17_port, QN => n56);
   position1_y_sum_reg_16_inst : DF3 port map( D => position1_n1594, C => 
                           CLK_top, Q => position1_y_sum_16_port, QN => n74);
   position1_y_sum_reg_15_inst : DF3 port map( D => position1_n1595, C => 
                           CLK_top, Q => position1_y_sum_15_port, QN => n57);
   position1_y_sum_reg_14_inst : DF3 port map( D => position1_n1596, C => 
                           CLK_top, Q => position1_y_sum_14_port, QN => n75);
   position1_y_sum_reg_13_inst : DF3 port map( D => position1_n1597, C => 
                           CLK_top, Q => position1_y_sum_13_port, QN => n58);
   position1_y_sum_reg_12_inst : DF3 port map( D => position1_n1598, C => 
                           CLK_top, Q => position1_y_sum_12_port, QN => n76);
   position1_y_sum_reg_11_inst : DF3 port map( D => position1_n1599, C => 
                           CLK_top, Q => position1_y_sum_11_port, QN => n59);
   position1_y_sum_reg_10_inst : DF3 port map( D => position1_n1600, C => 
                           CLK_top, Q => position1_y_sum_10_port, QN => n69);
   position1_y_sum_reg_9_inst : DF3 port map( D => position1_n1601, C => 
                           CLK_top, Q => position1_y_sum_9_port, QN => n51);
   position1_y_sum_reg_8_inst : DF3 port map( D => position1_n1602, C => 
                           CLK_top, Q => position1_y_sum_8_port, QN => n49);
   position1_y_sum_reg_7_inst : DF3 port map( D => position1_n1603, C => 
                           CLK_top, Q => position1_y_sum_7_port, QN => n93);
   position1_y_sum_reg_6_inst : DF3 port map( D => position1_n1604, C => 
                           CLK_top, Q => position1_y_sum_6_port, QN => n83);
   position1_y_sum_reg_5_inst : DF3 port map( D => position1_n1605, C => 
                           CLK_top, Q => position1_y_sum_5_port, QN => n84);
   position1_y_sum_reg_4_inst : DF3 port map( D => position1_n1606, C => 
                           CLK_top, Q => position1_y_sum_4_port, QN => n85);
   position1_y_sum_reg_3_inst : DF3 port map( D => position1_n1607, C => 
                           CLK_top, Q => position1_y_sum_3_port, QN => n94);
   position1_y_sum_reg_2_inst : DF3 port map( D => position1_n1608, C => 
                           CLK_top, Q => position1_y_sum_2_port, QN => n86);
   position1_y_sum_reg_1_inst : DF3 port map( D => position1_n1609, C => 
                           CLK_top, Q => position1_y_sum_1_port, QN => n87);
   position1_y_sum_reg_23_inst : DF3 port map( D => position1_n1587, C => 
                           CLK_top, Q => position1_y_sum_23_port, QN => n53);
   position1_y_sum_reg_24_inst : DF3 port map( D => position1_n1586, C => 
                           CLK_top, Q => position1_y_sum_24_port, QN => n99);
   position1_y_sum_reg_0_inst : DF3 port map( D => position1_n1610, C => 
                           CLK_top, Q => position1_N1938, QN => n97);
   position1_count_img_reg_19_inst : DF3 port map( D => n713, C => CLK_top, Q 
                           => position1_count_img_19_port, QN => n_1052);
   position1_count_img_reg_18_inst : DF3 port map( D => n712, C => CLK_top, Q 
                           => position1_count_img_18_port, QN => n_1053);
   position1_count_img_reg_17_inst : DF3 port map( D => n711, C => CLK_top, Q 
                           => position1_count_img_17_port, QN => n_1054);
   position1_count_img_reg_16_inst : DF3 port map( D => n710, C => CLK_top, Q 
                           => position1_count_img_16_port, QN => n_1055);
   position1_count_img_reg_15_inst : DF3 port map( D => n709, C => CLK_top, Q 
                           => position1_count_img_15_port, QN => n18);
   position1_count_img_reg_14_inst : DF3 port map( D => n708, C => CLK_top, Q 
                           => position1_count_img_14_port, QN => n_1056);
   position1_count_img_reg_13_inst : DF3 port map( D => n707, C => CLK_top, Q 
                           => position1_count_img_13_port, QN => n_1057);
   position1_count_img_reg_12_inst : DF3 port map( D => n706, C => CLK_top, Q 
                           => position1_count_img_12_port, QN => n_1058);
   position1_count_img_reg_11_inst : DF3 port map( D => n705, C => CLK_top, Q 
                           => position1_count_img_11_port, QN => n_1059);
   position1_count_img_reg_10_inst : DF3 port map( D => n704, C => CLK_top, Q 
                           => position1_count_img_10_port, QN => n_1060);
   position1_count_img_reg_9_inst : DF3 port map( D => n703, C => CLK_top, Q =>
                           position1_count_img_9_port, QN => n_1061);
   position1_count_img_reg_8_inst : DF3 port map( D => n702, C => CLK_top, Q =>
                           position1_count_img_8_port, QN => n_1062);
   position1_count_img_reg_7_inst : DF3 port map( D => n701, C => CLK_top, Q =>
                           position1_count_img_7_port, QN => n_1063);
   position1_count_img_reg_6_inst : DF3 port map( D => n700, C => CLK_top, Q =>
                           position1_count_img_6_port, QN => n_1064);
   position1_count_img_reg_5_inst : DF3 port map( D => n699, C => CLK_top, Q =>
                           position1_count_img_5_port, QN => n_1065);
   position1_count_img_reg_4_inst : DF3 port map( D => n698, C => CLK_top, Q =>
                           position1_count_img_4_port, QN => n_1066);
   position1_count_img_reg_3_inst : DF3 port map( D => n697, C => CLK_top, Q =>
                           position1_count_img_3_port, QN => n_1067);
   position1_count_img_reg_2_inst : DF3 port map( D => n696, C => CLK_top, Q =>
                           position1_count_img_2_port, QN => n_1068);
   position1_count_img_reg_1_inst : DF3 port map( D => n695, C => CLK_top, Q =>
                           position1_count_img_1_port, QN => n_1069);
   position1_state_reg_1_inst : DF3 port map( D => n486, C => CLK_top, Q => 
                           position1_state_1_port, QN => position1_n344);
   position1_state_reg_0_inst : DF3 port map( D => position1_N193, C => CLK_top
                           , Q => position1_state_0_port, QN => n_1070);
   position1_count_img_reg_0_inst : DF3 port map( D => n694, C => CLK_top, Q =>
                           position1_count_img_0_port, QN => position1_n802);
   position1_bi_reg_0_inst : DF3 port map( D => n725, C => CLK_top, Q => n_1071
                           , QN => position1_n370);
   position1_bi_reg_1_inst : DF3 port map( D => n724, C => CLK_top, Q => n_1072
                           , QN => position1_n369);
   position1_bi_reg_2_inst : DF3 port map( D => n723, C => CLK_top, Q => n_1073
                           , QN => position1_n368);
   position1_bi_reg_3_inst : DF3 port map( D => n722, C => CLK_top, Q => n_1074
                           , QN => position1_n367);
   position1_bi_reg_4_inst : DF3 port map( D => n721, C => CLK_top, Q => n_1075
                           , QN => position1_n366);
   position1_bi_reg_5_inst : DF3 port map( D => n720, C => CLK_top, Q => n_1076
                           , QN => position1_n365);
   position1_bi_reg_6_inst : DF3 port map( D => n719, C => CLK_top, Q => n_1077
                           , QN => position1_n364);
   position1_bi_reg_7_inst : DF3 port map( D => n718, C => CLK_top, Q => n_1078
                           , QN => position1_n363);
   position1_gi_reg_0_inst : DF3 port map( D => n733, C => CLK_top, Q => 
                           position1_gi_0_port, QN => position1_n362);
   position1_gi_reg_1_inst : DF3 port map( D => n732, C => CLK_top, Q => 
                           position1_gi_1_port, QN => n_1079);
   position1_gi_reg_2_inst : DF3 port map( D => n731, C => CLK_top, Q => 
                           position1_gi_2_port, QN => position1_n360);
   position1_gi_reg_3_inst : DF3 port map( D => n730, C => CLK_top, Q => 
                           position1_gi_3_port, QN => n_1080);
   position1_gi_reg_4_inst : DF3 port map( D => n729, C => CLK_top, Q => 
                           position1_gi_4_port, QN => position1_n358);
   position1_gi_reg_5_inst : DF3 port map( D => n728, C => CLK_top, Q => 
                           position1_gi_5_port, QN => position1_n357);
   position1_gi_reg_6_inst : DF3 port map( D => n727, C => CLK_top, Q => 
                           position1_gi_6_port, QN => position1_n356);
   position1_gi_reg_7_inst : DF3 port map( D => n726, C => CLK_top, Q => 
                           position1_gi_7_port, QN => n_1081);
   position1_ri_reg_0_inst : DF3 port map( D => n741, C => CLK_top, Q => n_1082
                           , QN => position1_n353);
   position1_ri_reg_1_inst : DF3 port map( D => n740, C => CLK_top, Q => n_1083
                           , QN => position1_n352);
   position1_ri_reg_2_inst : DF3 port map( D => n739, C => CLK_top, Q => n_1084
                           , QN => position1_n351);
   position1_ri_reg_3_inst : DF3 port map( D => n738, C => CLK_top, Q => n_1085
                           , QN => position1_n350);
   position1_ri_reg_4_inst : DF3 port map( D => n737, C => CLK_top, Q => n_1086
                           , QN => position1_n349);
   position1_ri_reg_5_inst : DF3 port map( D => n736, C => CLK_top, Q => n_1087
                           , QN => position1_n348);
   position1_ri_reg_6_inst : DF3 port map( D => n735, C => CLK_top, Q => n_1088
                           , QN => position1_n347);
   position1_ri_reg_7_inst : DF3 port map( D => n734, C => CLK_top, Q => n_1089
                           , QN => position1_n346);
   image_process1_r_out_reg_0_inst : DFE1 port map( D => image_process1_N8, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_0_port, 
                           QN => n_1090);
   image_process1_r_out_reg_1_inst : DFE1 port map( D => image_process1_N11, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_1_port, 
                           QN => n_1091);
   image_process1_r_out_reg_2_inst : DFE1 port map( D => image_process1_N14, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_2_port, 
                           QN => n_1092);
   image_process1_r_out_reg_3_inst : DFE1 port map( D => image_process1_N17, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_3_port, 
                           QN => n_1093);
   image_process1_r_out_reg_4_inst : DFE1 port map( D => image_process1_N20, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_4_port, 
                           QN => n_1094);
   image_process1_r_out_reg_5_inst : DFE1 port map( D => image_process1_N23, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_5_port, 
                           QN => n_1095);
   image_process1_r_out_reg_6_inst : DFE1 port map( D => image_process1_N26, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_6_port, 
                           QN => n_1096);
   image_process1_r_out_reg_7_inst : DFE1 port map( D => image_process1_N29, E 
                           => reset_top, C => CLK_top, Q => r_out_proc_7_port, 
                           QN => n_1097);
   image_process1_b_out_reg_0_inst : DFE1 port map( D => image_process1_N10, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_0_port, 
                           QN => n_1098);
   image_process1_b_out_reg_1_inst : DFE1 port map( D => 
                           image_process1_N13_port, E => reset_top, C => 
                           CLK_top, Q => b_out_proc_1_port, QN => n_1099);
   image_process1_b_out_reg_2_inst : DFE1 port map( D => image_process1_N16, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_2_port, 
                           QN => n_1100);
   image_process1_b_out_reg_3_inst : DFE1 port map( D => image_process1_N19, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_3_port, 
                           QN => n_1101);
   image_process1_b_out_reg_4_inst : DFE1 port map( D => image_process1_N22, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_4_port, 
                           QN => n_1102);
   image_process1_b_out_reg_5_inst : DFE1 port map( D => 
                           image_process1_N25_port, E => reset_top, C => 
                           CLK_top, Q => b_out_proc_5_port, QN => n_1103);
   image_process1_b_out_reg_6_inst : DFE1 port map( D => image_process1_N28, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_6_port, 
                           QN => n_1104);
   image_process1_b_out_reg_7_inst : DFE1 port map( D => image_process1_N31, E 
                           => reset_top, C => CLK_top, Q => b_out_proc_7_port, 
                           QN => n_1105);
   image_process1_g_out_reg_2_inst : DFE1 port map( D => n769, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_2_port, QN => n_1106);
   image_process1_g_out_reg_6_inst : DFE1 port map( D => n773, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_6_port, QN => n_1107);
   image_process1_g_out_reg_4_inst : DFE1 port map( D => n771, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_4_port, QN => n_1108);
   image_process1_g_out_reg_5_inst : DFE1 port map( D => n772, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_5_port, QN => n_1109);
   image_process1_g_out_reg_0_inst : DFE1 port map( D => n775, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_0_port, QN => n_1110);
   image_process1_g_out_reg_1_inst : DFE1 port map( D => n768, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_1_port, QN => n_1111);
   image_process1_g_out_reg_3_inst : DFE1 port map( D => n770, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_3_port, QN => n_1112);
   image_process1_g_out_reg_7_inst : DFE1 port map( D => n774, E => reset_top, 
                           C => CLK_top, Q => g_out_proc_7_port, QN => n_1113);
   position1_sub_226_U2_24 : XOR31 port map( A => position1_y_sum_24_port, B =>
                           n45, C => position1_sub_226_carry_24_port, Q => 
                           position1_N1962);
   position1_sub_216_U2_24 : XOR31 port map( A => position1_x_sum_24_port, B =>
                           n300, C => position1_sub_216_carry_24_port, Q => 
                           position1_N1545_port);
   position1_sub_226_I2_U2_24 : XOR31 port map( A => position1_N1987, B => n590
                           , C => position1_sub_226_I2_carry_24_port, Q => 
                           position1_N2014);
   position1_sub_216_I2_U2_24 : XOR31 port map( A => position1_N1570_port, B =>
                           n591, C => position1_sub_216_I2_carry_24_port, Q => 
                           position1_N1597_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_7 : MAJ31 port map( A => n491
                           , B => cam_x_7_port, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_7_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_8_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_3 : MAJ31 port map( A => n499
                           , B => cam_x_3_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_3_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_4_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_5 : MAJ31 port map( A => n495
                           , B => cam_x_5_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_5_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_6_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_1 : MAJ31 port map( A => n503
                           , B => cam_x_1_port, C => n505, Q => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_2_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_2 : MAJ31 port map( A => n501
                           , B => cam_x_2_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_2_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_3_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_5 : MAJ31 port map( A => n495
                           , B => cam_x_5_port, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_5_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_6_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_1 : MAJ31 port map( A => n503
                           , B => cam_x_1_port, C => cam_x_0_port, Q => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_2_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_3 : MAJ31 port map( A => 
                           cam_x_3_port, B => n499, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_3_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_4_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_2 : MAJ31 port map( A => 
                           cam_x_2_port, B => n501, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_2_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_3_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_6 : MAJ31 port map( A => n493
                           , B => cam_x_6_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_6_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_7_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_4 : MAJ31 port map( A => n497
                           , B => cam_x_4_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_4_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_5_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_6 : MAJ31 port map( A => n493
                           , B => cam_x_6_port, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_6_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_7_port);
   position1_dp_cluster_3_add_1_root_add_188_3_U1_4 : MAJ31 port map( A => n497
                           , B => cam_x_4_port, C => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_4_port, Q 
                           => 
                           position1_dp_cluster_3_add_1_root_add_188_3_carry_5_port);
   position1_dp_cluster_7_add_1_root_add_170_3_U1_7 : MAJ31 port map( A => n491
                           , B => cam_x_7_port, C => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_7_port, Q 
                           => 
                           position1_dp_cluster_7_add_1_root_add_170_3_carry_8_port);
   gensync1_comptY_reg_4_inst : DFE1 port map( D => gensync1_N60, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N169, QN 
                           => n13);
   gensync1_comptY_reg_3_inst : DFE1 port map( D => gensync1_N59, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N170, QN 
                           => n11);
   gensync1_comptY_reg_1_inst : DFE1 port map( D => gensync1_N57, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N172, QN 
                           => n9);
   gensync1_comptY_reg_2_inst : DFE1 port map( D => gensync1_N58, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N171, QN 
                           => n8);
   gensync1_comptY_reg_0_inst : DFE1 port map( D => gensync1_N56, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N173, QN 
                           => n3);
   gensync1_comptY_reg_5_inst : DFE1 port map( D => gensync1_N61, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N168, QN 
                           => n_1114);
   gensync1_comptY_reg_6_inst : DFE1 port map( D => gensync1_N62, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N167, QN 
                           => n_1115);
   gensync1_comptY_reg_7_inst : DFE1 port map( D => gensync1_N63, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N166, QN 
                           => n_1116);
   gensync1_comptY_reg_8_inst : DFE1 port map( D => gensync1_N64, E => 
                           gensync1_n107, C => CLK_top, Q => gensync1_N165, QN 
                           => n_1117);
   gensync1_comptY_reg_9_inst : DFE1 port map( D => gensync1_N65, E => 
                           gensync1_n107, C => CLK_top, Q => 
                           gensync1_comptY_9_port, QN => n_1118);
   U1 : XOR21 port map( A => position1_y_sum_9_port, B => 
                           position1_r409_carry_9_port, Q => 
                           position1_N364_port);
   U2 : XOR21 port map( A => position1_x_sum_9_port, B => 
                           position1_r406_carry_9_port, Q => position1_N289);
   U3 : NAND31 port map( A => position1_N267, B => IMG_top_port, C => 
                           position1_n1389, Q => position1_n1062);
   U4 : AOI221 port map( A => n1127, B => n549, C => position1_N1909, D => n553
                           , Q => position1_n1384);
   U5 : AOI221 port map( A => n908, B => n583, C => position1_N2326, D => n587,
                           Q => position1_n1208);
   U6 : NOR21 port map( A => gensync1_n102, B => n114, Q => gensync1_N31);
   U7 : NOR21 port map( A => n509, B => n113, Q => gensync1_N65);
   U8 : XOR21 port map( A => position1_x_sum_20_port, B => 
                           position1_r406_carry_20_port, Q => position1_N300);
   U9 : XOR21 port map( A => position1_x_sum_22_port, B => 
                           position1_r406_carry_22_port, Q => position1_N302);
   U10 : XOR21 port map( A => position1_x_sum_19_port, B => 
                           position1_r406_carry_19_port, Q => position1_N299);
   U11 : XOR21 port map( A => position1_x_sum_21_port, B => 
                           position1_r406_carry_21_port, Q => position1_N301);
   U12 : XOR21 port map( A => position1_x_sum_23_port, B => 
                           position1_r406_carry_23_port, Q => position1_N303);
   U13 : XOR21 port map( A => position1_x_sum_14_port, B => 
                           position1_r406_carry_14_port, Q => position1_N294);
   U14 : XOR21 port map( A => position1_x_sum_16_port, B => 
                           position1_r406_carry_16_port, Q => position1_N296);
   U15 : XOR21 port map( A => position1_x_sum_18_port, B => 
                           position1_r406_carry_18_port, Q => position1_N298);
   U16 : XOR21 port map( A => position1_y_sum_20_port, B => 
                           position1_r409_carry_20_port, Q => position1_N375);
   U17 : XOR21 port map( A => position1_y_sum_22_port, B => 
                           position1_r409_carry_22_port, Q => position1_N377);
   U18 : XOR21 port map( A => position1_x_sum_13_port, B => 
                           position1_r406_carry_13_port, Q => position1_N293);
   U19 : XOR21 port map( A => position1_x_sum_15_port, B => 
                           position1_r406_carry_15_port, Q => position1_N295);
   U20 : XOR21 port map( A => position1_x_sum_17_port, B => 
                           position1_r406_carry_17_port, Q => position1_N297);
   U21 : XOR21 port map( A => position1_y_sum_19_port, B => 
                           position1_r409_carry_19_port, Q => position1_N374);
   U22 : XOR21 port map( A => position1_y_sum_21_port, B => 
                           position1_r409_carry_21_port, Q => position1_N376);
   U23 : XOR21 port map( A => position1_y_sum_23_port, B => 
                           position1_r409_carry_23_port, Q => position1_N378);
   U24 : XOR21 port map( A => position1_x_sum_10_port, B => 
                           position1_r406_carry_10_port, Q => position1_N290);
   U25 : XOR21 port map( A => position1_x_sum_12_port, B => 
                           position1_r406_carry_12_port, Q => position1_N292);
   U26 : XOR21 port map( A => position1_y_sum_14_port, B => 
                           position1_r409_carry_14_port, Q => 
                           position1_N369_port);
   U27 : XOR21 port map( A => position1_y_sum_16_port, B => 
                           position1_r409_carry_16_port, Q => position1_N371);
   U28 : XOR21 port map( A => position1_y_sum_18_port, B => 
                           position1_r409_carry_18_port, Q => position1_N373);
   U29 : XOR21 port map( A => position1_y_sum_13_port, B => 
                           position1_r409_carry_13_port, Q => 
                           position1_N368_port);
   U30 : XOR21 port map( A => position1_y_sum_15_port, B => 
                           position1_r409_carry_15_port, Q => 
                           position1_N370_port);
   U31 : XOR21 port map( A => position1_y_sum_17_port, B => 
                           position1_r409_carry_17_port, Q => position1_N372);
   U32 : XOR21 port map( A => position1_x_sum_11_port, B => 
                           position1_r406_carry_11_port, Q => position1_N291);
   U33 : XOR21 port map( A => position1_y_sum_10_port, B => 
                           position1_r409_carry_10_port, Q => 
                           position1_N365_port);
   U34 : XOR21 port map( A => position1_y_sum_12_port, B => 
                           position1_r409_carry_12_port, Q => 
                           position1_N367_port);
   U35 : XOR21 port map( A => position1_y_sum_11_port, B => 
                           position1_r409_carry_11_port, Q => 
                           position1_N366_port);
   U36 : XOR21 port map( A => gensync1_N174, B => n477, Q => n34);
   U37 : OAI2111 port map( A => n2, B => n1712, C => n1048, D => 
                           position1_n1333, Q => position1_N2040);
   U38 : OAI2111 port map( A => n2, B => n2046, C => n1267, D => 
                           position1_n1529, Q => position1_N1623_port);
   U39 : INV3 port map( A => n103, Q => n1818);
   U40 : INV3 port map( A => n104, Q => n1484);
   U41 : INV3 port map( A => n109, Q => n2011);
   U42 : INV3 port map( A => n110, Q => n1677);
   U43 : INV3 port map( A => n111, Q => n2012);
   U44 : INV3 port map( A => n112, Q => n1678);
   U45 : BUF2 port map( A => n2128, Q => position1_dp_cluster_7_N314);
   U46 : BUF2 port map( A => position1_n1071, Q => n478);
   U47 : BUF2 port map( A => position1_N2457, Q => n469);
   U48 : BUF2 port map( A => position1_N2453, Q => n472);
   U49 : BUF2 port map( A => image_process1_n61, Q => n490);
   U50 : BUF2 port map( A => position1_N2449, Q => n475);
   U51 : BUF2 port map( A => position1_N2447, Q => n476);
   U52 : NOR40 port map( A => n1390, B => image_process1_gi_5_port, C => 
                           image_process1_gi_7_port, D => 
                           image_process1_gi_6_port, Q => 
                           image_process1_N59_port);
   U53 : NAND22 port map( A => gensync1_N9, B => n651, Q => gensync1_n102);
   U54 : BUF2 port map( A => position1_N194, Q => n486);
   U55 : INV3 port map( A => position1_n1500, Q => n1210);
   U56 : INV3 port map( A => position1_n1304, Q => n991);
   U57 : INV3 port map( A => position1_n1517, Q => n1228);
   U58 : INV3 port map( A => position1_n1321, Q => n1009);
   U59 : INV3 port map( A => position1_n1515, Q => n1226);
   U60 : INV3 port map( A => position1_n1319, Q => n1007);
   U61 : INV3 port map( A => position1_n1513, Q => n1224);
   U62 : INV3 port map( A => position1_n1317, Q => n1005);
   U63 : INV3 port map( A => position1_n1511, Q => n1222);
   U64 : INV3 port map( A => position1_n1315, Q => n1003);
   U65 : INV3 port map( A => position1_n1509, Q => n1220);
   U66 : INV3 port map( A => position1_n1313, Q => n1001);
   U67 : INV3 port map( A => position1_n1476, Q => n1183);
   U68 : INV3 port map( A => position1_n1280, Q => n964);
   U69 : INV3 port map( A => position1_n1519, Q => n1231);
   U70 : INV3 port map( A => position1_n1323, Q => n1012);
   U71 : INV3 port map( A => position1_n1443, Q => n1145);
   U72 : INV3 port map( A => position1_n1247, Q => n926);
   U73 : INV3 port map( A => position1_n1485, Q => n1194);
   U74 : INV3 port map( A => position1_n1289, Q => n975);
   U75 : INV3 port map( A => position1_n1469, Q => n1176);
   U76 : INV3 port map( A => position1_n1273, Q => n957);
   U77 : INV3 port map( A => position1_n1467, Q => n1174);
   U78 : INV3 port map( A => position1_n1271, Q => n955);
   U79 : INV3 port map( A => position1_n1465, Q => n1172);
   U80 : INV3 port map( A => position1_n1269, Q => n953);
   U81 : INV3 port map( A => position1_n1463, Q => n1170);
   U82 : INV3 port map( A => position1_n1267, Q => n951);
   U83 : INV3 port map( A => position1_n1461, Q => n1168);
   U84 : INV3 port map( A => position1_n1265, Q => n949);
   U85 : INV3 port map( A => position1_n1471, Q => n1178);
   U86 : INV3 port map( A => position1_n1275, Q => n959);
   U87 : INV3 port map( A => position1_n1495, Q => n1205);
   U88 : INV3 port map( A => position1_n1299, Q => n986);
   U89 : INV3 port map( A => position1_n1491, Q => n1201);
   U90 : INV3 port map( A => position1_n1295, Q => n982);
   U91 : INV3 port map( A => position1_n1489, Q => n1199);
   U92 : INV3 port map( A => position1_n1293, Q => n980);
   U93 : INV3 port map( A => position1_n1487, Q => n1197);
   U94 : INV3 port map( A => position1_n1291, Q => n978);
   U95 : INV3 port map( A => position1_n1445, Q => n1148);
   U96 : INV3 port map( A => position1_n1249, Q => n929);
   U97 : INV3 port map( A => position1_n1493, Q => n1203);
   U98 : INV3 port map( A => position1_n1297, Q => n984);
   U99 : NAND31 port map( A => position1_n1386, B => position1_n1384, C => 
                           position1_n1385, Q => n103);
   U100 : NAND31 port map( A => position1_n1210, B => position1_n1208, C => 
                           position1_n1209, Q => n104);
   U101 : NOR21 port map( A => position1_sub_216_I7_carry_23_port, B => n1162, 
                           Q => n125);
   U102 : NOR21 port map( A => position1_sub_226_I7_carry_23_port, B => n943, Q
                           => n141);
   U103 : NOR21 port map( A => position1_sub_216_I6_carry_23_port, B => n1188, 
                           Q => n121);
   U104 : NOR21 port map( A => position1_sub_226_I6_carry_23_port, B => n969, Q
                           => n137);
   U105 : INV3 port map( A => n124, Q => position1_sub_216_I7_carry_23_port);
   U106 : NOR21 port map( A => position1_sub_216_I7_carry_22_port, B => n1163, 
                           Q => n124);
   U107 : INV3 port map( A => n140, Q => position1_sub_226_I7_carry_23_port);
   U108 : NOR21 port map( A => position1_sub_226_I7_carry_22_port, B => n944, Q
                           => n140);
   U109 : INV3 port map( A => n128, Q => position1_sub_216_I8_carry_22_port);
   U110 : NOR21 port map( A => position1_sub_216_I8_carry_21_port, B => n1130, 
                           Q => n128);
   U111 : INV3 port map( A => n144, Q => position1_sub_226_I8_carry_22_port);
   U112 : NOR21 port map( A => position1_sub_226_I8_carry_21_port, B => n911, Q
                           => n144);
   U113 : INV3 port map( A => n129, Q => position1_sub_216_I8_carry_23_port);
   U114 : NOR21 port map( A => position1_sub_216_I8_carry_22_port, B => n1129, 
                           Q => n129);
   U115 : INV3 port map( A => n145, Q => position1_sub_226_I8_carry_23_port);
   U116 : NOR21 port map( A => position1_sub_226_I8_carry_22_port, B => n910, Q
                           => n145);
   U117 : INV3 port map( A => position1_n1421, Q => n1117);
   U118 : INV3 port map( A => position1_n1225, Q => n898);
   U119 : INV3 port map( A => position1_N2397, Q => n842);
   U120 : INV3 port map( A => position1_N2399, Q => n840);
   U121 : INV3 port map( A => position1_N2376, Q => n850);
   U122 : AOI221 port map( A => n535, B => position1_N1686, C => n533, D => 
                           position1_N1659, Q => position1_n1519);
   U123 : AOI221 port map( A => n569, B => position1_N2103, C => n567, D => 
                           position1_N2076, Q => position1_n1323);
   U124 : AOI221 port map( A => n547, B => position1_N1843, C => n545, D => 
                           n1175, Q => position1_n1443);
   U125 : AOI221 port map( A => n581, B => position1_N2260, C => n579, D => 
                           n956, Q => position1_n1247);
   U126 : AOI221 port map( A => n547, B => position1_N1841, C => n545, D => 
                           n1177, Q => position1_n1445);
   U127 : AOI221 port map( A => n581, B => position1_N2258, C => n579, D => 
                           n958, Q => position1_n1249);
   U128 : AOI221 port map( A => n540, B => position1_N1747, C => n537, D => 
                           n1221, Q => position1_n1485);
   U129 : AOI221 port map( A => n574, B => position1_N2164, C => n571, D => 
                           n1002, Q => position1_n1289);
   U130 : AOI221 port map( A => n1146, B => n549, C => position1_N1894, D => 
                           n551, Q => position1_n1419);
   U131 : AOI221 port map( A => n927, B => n583, C => position1_N2311, D => 
                           n585, Q => position1_n1223);
   U132 : AOI221 port map( A => n543, B => position1_N1790, C => n541, D => 
                           n1204, Q => position1_n1469);
   U133 : AOI221 port map( A => n577, B => position1_N2207, C => n575, D => 
                           n985, Q => position1_n1273);
   U134 : AOI221 port map( A => n543, B => position1_N1792, C => n541, D => 
                           n1202, Q => position1_n1467);
   U135 : AOI221 port map( A => n577, B => position1_N2209, C => n575, D => 
                           n983, Q => position1_n1271);
   U136 : AOI221 port map( A => n543, B => position1_N1794, C => n541, D => 
                           n1200, Q => position1_n1465);
   U137 : AOI221 port map( A => n577, B => position1_N2211, C => n575, D => 
                           n981, Q => position1_n1269);
   U138 : AOI221 port map( A => n544, B => position1_N1796, C => n541, D => 
                           n1198, Q => position1_n1463);
   U139 : AOI221 port map( A => n578, B => position1_N2213, C => n575, D => 
                           n979, Q => position1_n1267);
   U140 : AOI221 port map( A => n544, B => position1_N1798, C => n541, D => 
                           n1196, Q => position1_n1461);
   U141 : AOI221 port map( A => n578, B => position1_N2215, C => n575, D => 
                           n977, Q => position1_n1265);
   U142 : AOI221 port map( A => n543, B => position1_N1788, C => n541, D => 
                           n1206, Q => position1_n1471);
   U143 : AOI221 port map( A => n577, B => position1_N2205, C => n575, D => 
                           n987, Q => position1_n1275);
   U144 : AOI221 port map( A => n539, B => position1_N1737, C => n537, D => 
                           n1233, Q => position1_n1495);
   U145 : AOI221 port map( A => n573, B => position1_N2154, C => n571, D => 
                           n1014, Q => position1_n1299);
   U146 : AOI221 port map( A => n539, B => position1_N1741, C => n537, D => 
                           n1227, Q => position1_n1491);
   U147 : AOI221 port map( A => n573, B => position1_N2158, C => n571, D => 
                           n1008, Q => position1_n1295);
   U148 : AOI221 port map( A => n539, B => position1_N1743, C => n537, D => 
                           n1225, Q => position1_n1489);
   U149 : AOI221 port map( A => n573, B => position1_N2160, C => n571, D => 
                           n1006, Q => position1_n1293);
   U150 : AOI221 port map( A => n540, B => position1_N1745, C => n537, D => 
                           n1223, Q => position1_n1487);
   U151 : AOI221 port map( A => n574, B => position1_N2162, C => n571, D => 
                           n1004, Q => position1_n1291);
   U152 : AOI221 port map( A => n539, B => position1_N1739, C => n537, D => 
                           n1230, Q => position1_n1493);
   U153 : AOI221 port map( A => n573, B => position1_N2156, C => n571, D => 
                           n1011, Q => position1_n1297);
   U154 : AOI221 port map( A => n535, B => position1_N1688, C => n533, D => 
                           position1_N1661, Q => position1_n1517);
   U155 : AOI221 port map( A => n569, B => position1_N2105, C => n567, D => 
                           position1_N2078, Q => position1_n1321);
   U156 : AOI221 port map( A => n535, B => position1_N1690, C => n533, D => 
                           position1_N1663, Q => position1_n1515);
   U157 : AOI221 port map( A => n569, B => position1_N2107, C => n567, D => 
                           position1_N2080, Q => position1_n1319);
   U158 : AOI221 port map( A => n536, B => position1_N1692, C => n533, D => 
                           position1_N1665, Q => position1_n1513);
   U159 : AOI221 port map( A => n570, B => position1_N2109, C => n567, D => 
                           position1_N2082, Q => position1_n1317);
   U160 : AOI221 port map( A => n536, B => position1_N1694, C => n533, D => 
                           position1_N1667, Q => position1_n1511);
   U161 : AOI221 port map( A => n570, B => position1_N2111, C => n567, D => 
                           position1_N2084, Q => position1_n1315);
   U162 : AOI221 port map( A => n536, B => position1_N1696, C => n533, D => 
                           position1_N1669, Q => position1_n1509);
   U163 : AOI221 port map( A => n570, B => position1_N2113, C => n567, D => 
                           position1_N2086, Q => position1_n1313);
   U164 : AOI221 port map( A => n1144, B => n549, C => position1_N1896, D => 
                           n551, Q => position1_n1417);
   U165 : AOI221 port map( A => n925, B => n583, C => position1_N2313, D => 
                           n585, Q => position1_n1221);
   U166 : AOI221 port map( A => n1140, B => n549, C => position1_N1898, D => 
                           n552, Q => position1_n1415);
   U167 : AOI221 port map( A => n921, B => n583, C => position1_N2315, D => 
                           n586, Q => position1_n1219);
   U168 : AOI221 port map( A => n1137, B => n549, C => position1_N1900, D => 
                           n552, Q => position1_n1413);
   U169 : AOI221 port map( A => n918, B => n583, C => position1_N2317, D => 
                           n586, Q => position1_n1217);
   U170 : AOI221 port map( A => n538, B => n1242, C => n537, D => n1242, Q => 
                           position1_n1500);
   U171 : AOI221 port map( A => n572, B => n1023, C => n571, D => n1023, Q => 
                           position1_n1304);
   U172 : AOI221 port map( A => n1152, B => n549, C => position1_N1890, D => 
                           n551, Q => position1_n1423);
   U173 : AOI221 port map( A => n933, B => n583, C => position1_N2307, D => 
                           n585, Q => position1_n1227);
   U174 : AOI221 port map( A => n1149, B => n549, C => position1_N1892, D => 
                           n551, Q => position1_n1421);
   U175 : AOI221 port map( A => n930, B => n583, C => position1_N2309, D => 
                           n585, Q => position1_n1225);
   U176 : AOI221 port map( A => n542, B => n1211, C => n541, D => n1211, Q => 
                           position1_n1476);
   U177 : AOI221 port map( A => n576, B => n992, C => n575, D => n992, Q => 
                           position1_n1280);
   U178 : INV3 port map( A => n550, Q => n549);
   U179 : INV3 port map( A => n584, Q => n583);
   U180 : INV3 port map( A => n546, Q => n545);
   U181 : INV3 port map( A => n580, Q => n579);
   U182 : INV3 port map( A => n542, Q => n541);
   U183 : INV3 port map( A => n576, Q => n575);
   U184 : INV3 port map( A => n534, Q => n533);
   U185 : INV3 port map( A => n568, Q => n567);
   U186 : INV3 port map( A => n538, Q => n537);
   U187 : INV3 port map( A => n572, Q => n571);
   U188 : AOI221 port map( A => n1128, B => n549, C => position1_N1908, D => 
                           n553, Q => position1_n1385);
   U189 : XNR21 port map( A => n1128, B => position1_sub_216_I8_carry_23_port, 
                           Q => position1_N1908);
   U190 : XOR21 port map( A => n130, B => n1127, Q => position1_N1909);
   U191 : NOR21 port map( A => position1_sub_216_I8_carry_23_port, B => n1128, 
                           Q => n130);
   U192 : AOI221 port map( A => n1129, B => n549, C => position1_N1907, D => 
                           n553, Q => position1_n1386);
   U193 : XNR21 port map( A => n1129, B => position1_sub_216_I8_carry_22_port, 
                           Q => position1_N1907);
   U194 : AOI221 port map( A => n1130, B => n549, C => position1_N1906, D => 
                           n552, Q => position1_n1387);
   U195 : XNR21 port map( A => n1130, B => position1_sub_216_I8_carry_21_port, 
                           Q => position1_N1906);
   U196 : AOI221 port map( A => n909, B => n583, C => position1_N2325, D => 
                           n587, Q => position1_n1209);
   U197 : XNR21 port map( A => n909, B => position1_sub_226_I8_carry_23_port, Q
                           => position1_N2325);
   U198 : XOR21 port map( A => n146, B => n908, Q => position1_N2326);
   U199 : NOR21 port map( A => position1_sub_226_I8_carry_23_port, B => n909, Q
                           => n146);
   U200 : AOI221 port map( A => n910, B => n583, C => position1_N2324, D => 
                           n587, Q => position1_n1210);
   U201 : XNR21 port map( A => n910, B => position1_sub_226_I8_carry_22_port, Q
                           => position1_N2324);
   U202 : AOI221 port map( A => n911, B => n583, C => position1_N2323, D => 
                           n586, Q => position1_n1211);
   U203 : XNR21 port map( A => n911, B => position1_sub_226_I8_carry_21_port, Q
                           => position1_N2323);
   U204 : INV3 port map( A => position1_n1524, Q => n1241);
   U205 : INV3 port map( A => position1_n1328, Q => n1022);
   U206 : INV3 port map( A => position1_n1447, Q => n1151);
   U207 : AOI221 port map( A => n547, B => position1_N1839, C => n545, D => 
                           n1179, Q => position1_n1447);
   U208 : INV3 port map( A => position1_n1251, Q => n932);
   U209 : AOI221 port map( A => n581, B => position1_N2256, C => n579, D => 
                           n960, Q => position1_n1251);
   U210 : INV3 port map( A => position1_n1441, Q => n1142);
   U211 : AOI221 port map( A => n547, B => position1_N1845, C => n545, D => 
                           n1173, Q => position1_n1441);
   U212 : INV3 port map( A => position1_n1245, Q => n923);
   U213 : AOI221 port map( A => n581, B => position1_N2262, C => n579, D => 
                           n954, Q => position1_n1245);
   U214 : INV3 port map( A => position1_n1439, Q => n1139);
   U215 : AOI221 port map( A => n547, B => position1_N1847, C => n545, D => 
                           n1171, Q => position1_n1439);
   U216 : INV3 port map( A => position1_n1243, Q => n920);
   U217 : AOI221 port map( A => n581, B => position1_N2264, C => n579, D => 
                           n952, Q => position1_n1243);
   U218 : INV3 port map( A => position1_n1437, Q => n1136);
   U219 : AOI221 port map( A => n548, B => position1_N1849, C => n545, D => 
                           n1169, Q => position1_n1437);
   U220 : INV3 port map( A => position1_n1241, Q => n917);
   U221 : AOI221 port map( A => n582, B => position1_N2266, C => n579, D => 
                           n950, Q => position1_n1241);
   U222 : INV3 port map( A => n530, Q => n528);
   U223 : INV3 port map( A => n564, Q => n562);
   U224 : INV3 port map( A => position1_n1516, Q => n1227);
   U225 : INV3 port map( A => position1_n1320, Q => n1008);
   U226 : INV3 port map( A => position1_n1514, Q => n1225);
   U227 : INV3 port map( A => position1_n1318, Q => n1006);
   U228 : INV3 port map( A => position1_n1512, Q => n1223);
   U229 : INV3 port map( A => position1_n1316, Q => n1004);
   U230 : INV3 port map( A => position1_n1510, Q => n1221);
   U231 : INV3 port map( A => position1_n1314, Q => n1002);
   U232 : INV3 port map( A => position1_n1508, Q => n1219);
   U233 : INV3 port map( A => position1_n1312, Q => n1000);
   U234 : INV3 port map( A => position1_n1456, Q => n1163);
   U235 : AOI221 port map( A => n544, B => position1_N1803, C => n541, D => 
                           n1189, Q => position1_n1456);
   U236 : XNR21 port map( A => n1189, B => position1_sub_216_I6_carry_22_port, 
                           Q => position1_N1803);
   U237 : INV3 port map( A => position1_n1260, Q => n944);
   U238 : AOI221 port map( A => n578, B => position1_N2220, C => n575, D => 
                           n970, Q => position1_n1260);
   U239 : XNR21 port map( A => n970, B => position1_sub_226_I6_carry_22_port, Q
                           => position1_N2220);
   U240 : INV3 port map( A => position1_n1455, Q => n1162);
   U241 : AOI221 port map( A => n544, B => position1_N1804, C => n541, D => 
                           n1188, Q => position1_n1455);
   U242 : XNR21 port map( A => n1188, B => position1_sub_216_I6_carry_23_port, 
                           Q => position1_N1804);
   U243 : INV3 port map( A => position1_n1259, Q => n943);
   U244 : AOI221 port map( A => n578, B => position1_N2221, C => n575, D => 
                           n969, Q => position1_n1259);
   U245 : XNR21 port map( A => n969, B => position1_sub_226_I6_carry_23_port, Q
                           => position1_N2221);
   U246 : INV3 port map( A => position1_n1460, Q => n1167);
   U247 : INV3 port map( A => position1_n1264, Q => n948);
   U248 : INV3 port map( A => position1_n1494, Q => n1204);
   U249 : INV3 port map( A => position1_n1298, Q => n985);
   U250 : INV3 port map( A => position1_n1492, Q => n1202);
   U251 : INV3 port map( A => position1_n1296, Q => n983);
   U252 : INV3 port map( A => position1_n1490, Q => n1200);
   U253 : INV3 port map( A => position1_n1294, Q => n981);
   U254 : INV3 port map( A => position1_n1488, Q => n1198);
   U255 : INV3 port map( A => position1_n1292, Q => n979);
   U256 : INV3 port map( A => position1_n1486, Q => n1196);
   U257 : INV3 port map( A => position1_n1290, Q => n977);
   U258 : INV3 port map( A => position1_n1498, Q => n1208);
   U259 : INV3 port map( A => position1_n1302, Q => n989);
   U260 : INV3 port map( A => position1_n1496, Q => n1206);
   U261 : INV3 port map( A => position1_n1300, Q => n987);
   U262 : INV3 port map( A => position1_n1432, Q => n1130);
   U263 : AOI221 port map( A => n548, B => position1_N1854, C => n545, D => 
                           n1164, Q => position1_n1432);
   U264 : XNR21 port map( A => n1164, B => position1_sub_216_I7_carry_21_port, 
                           Q => position1_N1854);
   U265 : INV3 port map( A => position1_n1431, Q => n1129);
   U266 : AOI221 port map( A => n548, B => position1_N1855, C => n545, D => 
                           n1163, Q => position1_n1431);
   U267 : XNR21 port map( A => n1163, B => position1_sub_216_I7_carry_22_port, 
                           Q => position1_N1855);
   U268 : INV3 port map( A => position1_n1236, Q => n911);
   U269 : AOI221 port map( A => n582, B => position1_N2271, C => n579, D => 
                           n945, Q => position1_n1236);
   U270 : XNR21 port map( A => n945, B => position1_sub_226_I7_carry_21_port, Q
                           => position1_N2271);
   U271 : INV3 port map( A => position1_n1235, Q => n910);
   U272 : AOI221 port map( A => n582, B => position1_N2272, C => n579, D => 
                           n944, Q => position1_n1235);
   U273 : XNR21 port map( A => n944, B => position1_sub_226_I7_carry_22_port, Q
                           => position1_N2272);
   U274 : INV3 port map( A => position1_n1430, Q => n1128);
   U275 : AOI221 port map( A => n548, B => position1_N1856, C => n545, D => 
                           n1162, Q => position1_n1430);
   U276 : XNR21 port map( A => n1162, B => position1_sub_216_I7_carry_23_port, 
                           Q => position1_N1856);
   U277 : INV3 port map( A => position1_n1234, Q => n909);
   U278 : AOI221 port map( A => n582, B => position1_N2273, C => n579, D => 
                           n943, Q => position1_n1234);
   U279 : XNR21 port map( A => n943, B => position1_sub_226_I7_carry_23_port, Q
                           => position1_N2273);
   U280 : INV3 port map( A => position1_n1459, Q => n1166);
   U281 : INV3 port map( A => position1_n1263, Q => n947);
   U282 : INV3 port map( A => position1_n1520, Q => n1233);
   U283 : INV3 port map( A => position1_n1324, Q => n1014);
   U284 : INV3 port map( A => position1_n1473, Q => n1180);
   U285 : INV3 port map( A => position1_n1277, Q => n961);
   U286 : INV3 port map( A => position1_n1480, Q => n1188);
   U287 : AOI221 port map( A => n540, B => position1_N1752, C => n537, D => 
                           n1216, Q => position1_n1480);
   U288 : XNR21 port map( A => n1216, B => position1_sub_216_I5_carry_23_port, 
                           Q => position1_N1752);
   U289 : INV3 port map( A => position1_n1284, Q => n969);
   U290 : AOI221 port map( A => n574, B => position1_N2169, C => n571, D => 
                           n997, Q => position1_n1284);
   U291 : XNR21 port map( A => n997, B => position1_sub_226_I5_carry_23_port, Q
                           => position1_N2169);
   U292 : INV3 port map( A => position1_n1522, Q => n1237);
   U293 : INV3 port map( A => position1_n1326, Q => n1018);
   U294 : INV3 port map( A => position1_n1435, Q => n1134);
   U295 : INV3 port map( A => position1_n1239, Q => n915);
   U296 : INV3 port map( A => position1_n1497, Q => n1207);
   U297 : INV3 port map( A => position1_n1301, Q => n988);
   U298 : INV3 port map( A => n530, Q => n529);
   U299 : INV3 port map( A => n564, Q => n563);
   U300 : INV3 port map( A => position1_n1452, Q => n1159);
   U301 : AOI221 port map( A => n546, B => n1184, C => n545, D => n1184, Q => 
                           position1_n1452);
   U302 : INV3 port map( A => position1_n1256, Q => n940);
   U303 : AOI221 port map( A => n580, B => n965, C => n579, D => n965, Q => 
                           position1_n1256);
   U304 : INV3 port map( A => position1_n1436, Q => n1135);
   U305 : INV3 port map( A => position1_n1240, Q => n916);
   U306 : INV3 port map( A => position1_n1474, Q => n1181);
   U307 : INV3 port map( A => position1_n1278, Q => n962);
   U308 : INV3 port map( A => position1_n1472, Q => n1179);
   U309 : INV3 port map( A => position1_n1276, Q => n960);
   U310 : INV3 port map( A => position1_n1470, Q => n1177);
   U311 : INV3 port map( A => position1_n1274, Q => n958);
   U312 : INV3 port map( A => position1_n1466, Q => n1173);
   U313 : INV3 port map( A => position1_n1270, Q => n954);
   U314 : INV3 port map( A => position1_n1464, Q => n1171);
   U315 : INV3 port map( A => position1_n1268, Q => n952);
   U316 : INV3 port map( A => position1_n1462, Q => n1169);
   U317 : INV3 port map( A => position1_n1266, Q => n950);
   U318 : INV3 port map( A => position1_n1468, Q => n1175);
   U319 : INV3 port map( A => position1_n1272, Q => n956);
   U320 : INV3 port map( A => position1_n1507, Q => n1218);
   U321 : INV3 port map( A => position1_n1311, Q => n999);
   U322 : INV3 port map( A => position1_n1450, Q => n1155);
   U323 : INV3 port map( A => position1_n1254, Q => n936);
   U324 : INV3 port map( A => position1_n1448, Q => n1152);
   U325 : INV3 port map( A => position1_n1252, Q => n933);
   U326 : INV3 port map( A => position1_n1446, Q => n1149);
   U327 : INV3 port map( A => position1_n1250, Q => n930);
   U328 : INV3 port map( A => position1_n1440, Q => n1140);
   U329 : INV3 port map( A => position1_n1244, Q => n921);
   U330 : INV3 port map( A => position1_n1438, Q => n1137);
   U331 : INV3 port map( A => position1_n1242, Q => n918);
   U332 : INV3 port map( A => position1_n1454, Q => n1161);
   U333 : AOI221 port map( A => n544, B => position1_N1805, C => n541, D => 
                           n1187, Q => position1_n1454);
   U334 : XNR21 port map( A => position1_sub_216_I6_carry_24_port, B => n1187, 
                           Q => position1_N1805);
   U335 : INV3 port map( A => n121, Q => position1_sub_216_I6_carry_24_port);
   U336 : INV3 port map( A => position1_n1258, Q => n942);
   U337 : AOI221 port map( A => n578, B => position1_N2222, C => n575, D => 
                           n968, Q => position1_n1258);
   U338 : XNR21 port map( A => position1_sub_226_I6_carry_24_port, B => n968, Q
                           => position1_N2222);
   U339 : INV3 port map( A => n137, Q => position1_sub_226_I6_carry_24_port);
   U340 : INV3 port map( A => position1_n1429, Q => n1127);
   U341 : AOI221 port map( A => n548, B => position1_N1857, C => n545, D => 
                           n1161, Q => position1_n1429);
   U342 : XNR21 port map( A => position1_sub_216_I7_carry_24_port, B => n1161, 
                           Q => position1_N1857);
   U343 : INV3 port map( A => n125, Q => position1_sub_216_I7_carry_24_port);
   U344 : INV3 port map( A => position1_n1233, Q => n908);
   U345 : AOI221 port map( A => n582, B => position1_N2274, C => n579, D => 
                           n942, Q => position1_n1233);
   U346 : XNR21 port map( A => position1_sub_226_I7_carry_24_port, B => n942, Q
                           => position1_N2274);
   U347 : INV3 port map( A => n141, Q => position1_sub_226_I7_carry_24_port);
   U348 : INV3 port map( A => position1_n1479, Q => n1187);
   U349 : AOI221 port map( A => n540, B => position1_N1753, C => n537, D => 
                           n1215, Q => position1_n1479);
   U350 : XNR21 port map( A => position1_sub_216_I5_carry_24_port, B => n1215, 
                           Q => position1_N1753);
   U351 : INV3 port map( A => n118, Q => position1_sub_216_I5_carry_24_port);
   U352 : INV3 port map( A => position1_n1283, Q => n968);
   U353 : AOI221 port map( A => n574, B => position1_N2170, C => n571, D => 
                           n996, Q => position1_n1283);
   U354 : XNR21 port map( A => position1_sub_226_I5_carry_24_port, B => n996, Q
                           => position1_N2170);
   U355 : INV3 port map( A => n134, Q => position1_sub_226_I5_carry_24_port);
   U356 : INV3 port map( A => position1_n1453, Q => n1160);
   U357 : AOI221 port map( A => n546, B => n1185, C => n545, D => n1185, Q => 
                           position1_n1453);
   U358 : INV3 port map( A => position1_n1257, Q => n941);
   U359 : AOI221 port map( A => n580, B => n966, C => n579, D => n966, Q => 
                           position1_n1257);
   U360 : INV3 port map( A => position1_n1502, Q => n1212);
   U361 : AOI221 port map( A => n538, B => n1244, C => n537, D => n1244, Q => 
                           position1_n1502);
   U362 : INV3 port map( A => position1_n1501, Q => n1211);
   U363 : AOI221 port map( A => n538, B => n1243, C => n537, D => n1243, Q => 
                           position1_n1501);
   U364 : INV3 port map( A => position1_n1503, Q => n1213);
   U365 : AOI221 port map( A => n538, B => n1245, C => n537, D => n1245, Q => 
                           position1_n1503);
   U366 : INV3 port map( A => position1_n1306, Q => n993);
   U367 : AOI221 port map( A => n572, B => n1025, C => n571, D => n1025, Q => 
                           position1_n1306);
   U368 : INV3 port map( A => position1_n1305, Q => n992);
   U369 : AOI221 port map( A => n572, B => n1024, C => n571, D => n1024, Q => 
                           position1_n1305);
   U370 : INV3 port map( A => position1_n1307, Q => n994);
   U371 : AOI221 port map( A => n572, B => n1026, C => n571, D => n1026, Q => 
                           position1_n1307);
   U372 : INV3 port map( A => position1_n1478, Q => n1185);
   U373 : AOI221 port map( A => n542, B => n1213, C => n541, D => n1213, Q => 
                           position1_n1478);
   U374 : INV3 port map( A => position1_n1477, Q => n1184);
   U375 : AOI221 port map( A => n542, B => n1212, C => n541, D => n1212, Q => 
                           position1_n1477);
   U376 : INV3 port map( A => position1_n1282, Q => n966);
   U377 : AOI221 port map( A => n576, B => n994, C => n575, D => n994, Q => 
                           position1_n1282);
   U378 : INV3 port map( A => position1_n1281, Q => n965);
   U379 : AOI221 port map( A => n576, B => n993, C => n575, D => n993, Q => 
                           position1_n1281);
   U380 : NOR21 port map( A => position1_sub_216_I5_carry_23_port, B => n1216, 
                           Q => n118);
   U381 : NOR21 port map( A => position1_sub_226_I5_carry_23_port, B => n997, Q
                           => n134);
   U382 : XNR21 port map( A => n1131, B => position1_sub_216_I8_carry_20_port, 
                           Q => position1_N1905);
   U383 : XNR21 port map( A => n912, B => position1_sub_226_I8_carry_20_port, Q
                           => position1_N2322);
   U384 : BUF2 port map( A => n532, Q => n531);
   U385 : BUF2 port map( A => n566, Q => n565);
   U386 : INV3 port map( A => n120, Q => position1_sub_216_I6_carry_23_port);
   U387 : NOR21 port map( A => position1_sub_216_I6_carry_22_port, B => n1189, 
                           Q => n120);
   U388 : INV3 port map( A => n136, Q => position1_sub_226_I6_carry_23_port);
   U389 : NOR21 port map( A => position1_sub_226_I6_carry_22_port, B => n970, Q
                           => n136);
   U390 : INV3 port map( A => n123, Q => position1_sub_216_I7_carry_22_port);
   U391 : NOR21 port map( A => position1_sub_216_I7_carry_21_port, B => n1164, 
                           Q => n123);
   U392 : INV3 port map( A => n127, Q => position1_sub_216_I8_carry_21_port);
   U393 : NOR21 port map( A => position1_sub_216_I8_carry_20_port, B => n1131, 
                           Q => n127);
   U394 : INV3 port map( A => n139, Q => position1_sub_226_I7_carry_22_port);
   U395 : NOR21 port map( A => position1_sub_226_I7_carry_21_port, B => n945, Q
                           => n139);
   U396 : INV3 port map( A => n143, Q => position1_sub_226_I8_carry_21_port);
   U397 : NOR21 port map( A => position1_sub_226_I8_carry_20_port, B => n912, Q
                           => n143);
   U398 : INV3 port map( A => position1_n1416, Q => n1111);
   U399 : INV3 port map( A => position1_n1220, Q => n892);
   U400 : INV3 port map( A => position1_n1414, Q => n1109);
   U401 : INV3 port map( A => position1_n1218, Q => n890);
   U402 : INV3 port map( A => position1_n1426, Q => n1122);
   U403 : INV3 port map( A => position1_n1230, Q => n903);
   U404 : INV3 port map( A => position1_n1424, Q => n1120);
   U405 : INV3 port map( A => position1_n1228, Q => n901);
   U406 : INV3 port map( A => position1_n1422, Q => n1118);
   U407 : INV3 port map( A => position1_n1226, Q => n899);
   U408 : NOR21 port map( A => n1103, B => n1104, Q => n1819);
   U409 : INV3 port map( A => position1_n1388, Q => n1104);
   U410 : INV3 port map( A => position1_n1387, Q => n1103);
   U411 : AOI221 port map( A => n1131, B => n549, C => position1_N1905, D => 
                           n552, Q => position1_n1388);
   U412 : NOR21 port map( A => n884, B => n885, Q => n1485);
   U413 : INV3 port map( A => position1_n1212, Q => n885);
   U414 : INV3 port map( A => position1_n1211, Q => n884);
   U415 : AOI221 port map( A => n912, B => n583, C => position1_N2322, D => 
                           n586, Q => position1_n1212);
   U416 : INV3 port map( A => position1_n1428, Q => n1124);
   U417 : AOI221 port map( A => n1160, B => n549, C => n1160, D => n550, Q => 
                           position1_n1428);
   U418 : INV3 port map( A => position1_n1232, Q => n905);
   U419 : AOI221 port map( A => n941, B => n583, C => n941, D => n584, Q => 
                           position1_n1232);
   U420 : XOR21 port map( A => n497, B => position1_add_250_carry_4_port, Q => 
                           position1_N2397);
   U421 : XOR21 port map( A => n493, B => position1_add_250_carry_6_port, Q => 
                           position1_N2399);
   U422 : XNR21 port map( A => n497, B => position1_sub_250_carry_4_port, Q => 
                           position1_N2376);
   U423 : XNR21 port map( A => n493, B => position1_sub_250_carry_6_port, Q => 
                           position1_N2378);
   U424 : BUF2 port map( A => position1_n856, Q => n639);
   U425 : BUF2 port map( A => position1_n856, Q => n638);
   U426 : BUF2 port map( A => position1_n856, Q => n637);
   U427 : NAND22 port map( A => n743, B => n784, Q => position1_n1057);
   U428 : BUF2 port map( A => n742, Q => n513);
   U429 : NOR21 port map( A => n311, B => n312, Q => 
                           position1_add_250_carry_7_port);
   U430 : INV3 port map( A => n493, Q => n312);
   U431 : INV3 port map( A => position1_add_250_carry_6_port, Q => n311);
   U432 : BUF2 port map( A => n742, Q => n514);
   U433 : INV3 port map( A => n151, Q => position1_sub_250_carry_7_port);
   U434 : NOR21 port map( A => position1_sub_250_carry_6_port, B => n493, Q => 
                           n151);
   U435 : INV3 port map( A => n149, Q => position1_sub_250_carry_5_port);
   U436 : NOR21 port map( A => position1_sub_250_carry_4_port, B => n497, Q => 
                           n149);
   U437 : INV3 port map( A => position1_N2401, Q => n838);
   U438 : INV3 port map( A => position1_N2409, Q => n795);
   U439 : INV3 port map( A => position1_N2398, Q => n841);
   U440 : INV3 port map( A => position1_N2400, Q => n839);
   U441 : INV3 port map( A => position1_N2380, Q => n846);
   U442 : INV3 port map( A => position1_N2377, Q => n849);
   U443 : INV3 port map( A => position1_N2379, Q => n847);
   U444 : NOR21 port map( A => n307, B => n308, Q => 
                           position1_add_250_carry_5_port);
   U445 : INV3 port map( A => n497, Q => n308);
   U446 : INV3 port map( A => position1_add_250_carry_4_port, Q => n307);
   U447 : BUF2 port map( A => position1_n859, Q => n647);
   U448 : BUF2 port map( A => position1_n859, Q => n648);
   U449 : BUF2 port map( A => position1_n859, Q => n649);
   U450 : BUF2 port map( A => position1_n856, Q => n640);
   U451 : INV3 port map( A => image_process1_n97, Q => n778);
   U452 : INV3 port map( A => position1_N1634_port, Q => n1294);
   U453 : INV3 port map( A => position1_N2051, Q => n1075);
   U454 : INV3 port map( A => position1_N1636, Q => n1289);
   U455 : INV3 port map( A => position1_N2053, Q => n1070);
   U456 : INV3 port map( A => position1_N1638, Q => n1285);
   U457 : INV3 port map( A => position1_N2055, Q => n1066);
   U458 : INV3 port map( A => position1_N1640, Q => n1281);
   U459 : INV3 port map( A => position1_N2057, Q => n1062);
   U460 : INV3 port map( A => position1_N1642, Q => n1277);
   U461 : INV3 port map( A => position1_N2059, Q => n1058);
   U462 : INV3 port map( A => position1_N1644, Q => n1273);
   U463 : INV3 port map( A => position1_N2061, Q => n1054);
   U464 : INV3 port map( A => position1_N1646, Q => n1250);
   U465 : INV3 port map( A => position1_N2063, Q => n1031);
   U466 : INV3 port map( A => position1_N1648, Q => n1247);
   U467 : INV3 port map( A => position1_N2065, Q => n1028);
   U468 : AOI221 port map( A => n544, B => position1_N1799, C => n541, D => 
                           n1194, Q => position1_n1460);
   U469 : AOI221 port map( A => n578, B => position1_N2216, C => n575, D => 
                           n975, Q => position1_n1264);
   U470 : AOI221 port map( A => n548, B => position1_N1851, C => n545, D => 
                           n1167, Q => position1_n1435);
   U471 : AOI221 port map( A => n582, B => position1_N2268, C => n579, D => 
                           n948, Q => position1_n1239);
   U472 : AOI221 port map( A => n544, B => position1_N1800, C => n541, D => 
                           n1193, Q => position1_n1459);
   U473 : AOI221 port map( A => n578, B => position1_N2217, C => n575, D => 
                           n974, Q => position1_n1263);
   U474 : AOI221 port map( A => n535, B => position1_N1685, C => n533, D => 
                           position1_N1658, Q => position1_n1520);
   U475 : AOI221 port map( A => n569, B => position1_N2102, C => n567, D => 
                           position1_N2075, Q => position1_n1324);
   U476 : AOI221 port map( A => n535, B => position1_N1683, C => n533, D => 
                           position1_N1656, Q => position1_n1522);
   U477 : AOI221 port map( A => n569, B => position1_N2100, C => n567, D => 
                           position1_N2073, Q => position1_n1326);
   U478 : AOI221 port map( A => n548, B => position1_N1850, C => n545, D => 
                           n1168, Q => position1_n1436);
   U479 : AOI221 port map( A => n582, B => position1_N2267, C => n579, D => 
                           n949, Q => position1_n1240);
   U480 : AOI221 port map( A => n535, B => position1_N1654, C => n533, D => 
                           position1_N1654, Q => position1_n1524);
   U481 : AOI221 port map( A => n569, B => position1_N2071, C => n567, D => 
                           position1_N2071, Q => position1_n1328);
   U482 : AOI221 port map( A => n543, B => position1_N1786, C => n541, D => 
                           n1208, Q => position1_n1473);
   U483 : AOI221 port map( A => n577, B => position1_N2203, C => n575, D => 
                           n989, Q => position1_n1277);
   U484 : AOI221 port map( A => n539, B => position1_N1735, C => n537, D => 
                           n1237, Q => position1_n1497);
   U485 : AOI221 port map( A => n573, B => position1_N2152, C => n571, D => 
                           n1018, Q => position1_n1301);
   U486 : AOI221 port map( A => n1142, B => n549, C => position1_N1897, D => 
                           n551, Q => position1_n1416);
   U487 : AOI221 port map( A => n923, B => n583, C => position1_N2314, D => 
                           n585, Q => position1_n1220);
   U488 : AOI221 port map( A => n1139, B => n549, C => position1_N1899, D => 
                           n552, Q => position1_n1414);
   U489 : AOI221 port map( A => n920, B => n583, C => position1_N2316, D => 
                           n586, Q => position1_n1218);
   U490 : AOI221 port map( A => n1136, B => n549, C => position1_N1901, D => 
                           n552, Q => position1_n1412);
   U491 : AOI221 port map( A => n917, B => n583, C => position1_N2318, D => 
                           n586, Q => position1_n1216);
   U492 : AOI221 port map( A => n1157, B => n549, C => position1_N1887, D => 
                           n550, Q => position1_n1426);
   U493 : AOI221 port map( A => n938, B => n583, C => position1_N2304, D => 
                           n584, Q => position1_n1230);
   U494 : AOI221 port map( A => n1154, B => n549, C => position1_N1889, D => 
                           n551, Q => position1_n1424);
   U495 : AOI221 port map( A => n935, B => n583, C => position1_N2306, D => 
                           n585, Q => position1_n1228);
   U496 : AOI221 port map( A => n1151, B => n549, C => position1_N1891, D => 
                           n551, Q => position1_n1422);
   U497 : AOI221 port map( A => n932, B => n583, C => position1_N2308, D => 
                           n585, Q => position1_n1226);
   U498 : AOI221 port map( A => n536, B => position1_N1698, C => n533, D => 
                           position1_N1671, Q => position1_n1507);
   U499 : AOI221 port map( A => n570, B => position1_N2115, C => n567, D => 
                           position1_N2088, Q => position1_n1311);
   U500 : AOI221 port map( A => n535, B => position1_N1689, C => n533, D => 
                           position1_N1662, Q => position1_n1516);
   U501 : AOI221 port map( A => n569, B => position1_N2106, C => n567, D => 
                           position1_N2079, Q => position1_n1320);
   U502 : AOI221 port map( A => n535, B => position1_N1691, C => n533, D => 
                           position1_N1664, Q => position1_n1514);
   U503 : AOI221 port map( A => n569, B => position1_N2108, C => n567, D => 
                           position1_N2081, Q => position1_n1318);
   U504 : AOI221 port map( A => n536, B => position1_N1693, C => n533, D => 
                           position1_N1666, Q => position1_n1512);
   U505 : AOI221 port map( A => n570, B => position1_N2110, C => n567, D => 
                           position1_N2083, Q => position1_n1316);
   U506 : AOI221 port map( A => n536, B => position1_N1695, C => n533, D => 
                           position1_N1668, Q => position1_n1510);
   U507 : AOI221 port map( A => n570, B => position1_N2112, C => n567, D => 
                           position1_N2085, Q => position1_n1314);
   U508 : AOI221 port map( A => n536, B => position1_N1697, C => n533, D => 
                           position1_N1670, Q => position1_n1508);
   U509 : AOI221 port map( A => n570, B => position1_N2114, C => n567, D => 
                           position1_N2087, Q => position1_n1312);
   U510 : AOI221 port map( A => n543, B => position1_N1785, C => n541, D => 
                           n1209, Q => position1_n1474);
   U511 : AOI221 port map( A => n577, B => position1_N2202, C => n575, D => 
                           n990, Q => position1_n1278);
   U512 : AOI221 port map( A => n543, B => position1_N1787, C => n541, D => 
                           n1207, Q => position1_n1472);
   U513 : AOI221 port map( A => n577, B => position1_N2204, C => n575, D => 
                           n988, Q => position1_n1276);
   U514 : AOI221 port map( A => n543, B => position1_N1789, C => n541, D => 
                           n1205, Q => position1_n1470);
   U515 : AOI221 port map( A => n577, B => position1_N2206, C => n575, D => 
                           n986, Q => position1_n1274);
   U516 : AOI221 port map( A => n543, B => position1_N1793, C => n541, D => 
                           n1201, Q => position1_n1466);
   U517 : AOI221 port map( A => n577, B => position1_N2210, C => n575, D => 
                           n982, Q => position1_n1270);
   U518 : AOI221 port map( A => n543, B => position1_N1795, C => n541, D => 
                           n1199, Q => position1_n1464);
   U519 : AOI221 port map( A => n577, B => position1_N2212, C => n575, D => 
                           n980, Q => position1_n1268);
   U520 : AOI221 port map( A => n544, B => position1_N1797, C => n541, D => 
                           n1197, Q => position1_n1462);
   U521 : AOI221 port map( A => n578, B => position1_N2214, C => n575, D => 
                           n978, Q => position1_n1266);
   U522 : AOI221 port map( A => n543, B => position1_N1791, C => n541, D => 
                           n1203, Q => position1_n1468);
   U523 : AOI221 port map( A => n577, B => position1_N2208, C => n575, D => 
                           n984, Q => position1_n1272);
   U524 : AOI221 port map( A => n539, B => position1_N1738, C => n537, D => 
                           n1231, Q => position1_n1494);
   U525 : AOI221 port map( A => n573, B => position1_N2155, C => n571, D => 
                           n1012, Q => position1_n1298);
   U526 : AOI221 port map( A => n539, B => position1_N1740, C => n537, D => 
                           n1228, Q => position1_n1492);
   U527 : AOI221 port map( A => n573, B => position1_N2157, C => n571, D => 
                           n1009, Q => position1_n1296);
   U528 : AOI221 port map( A => n539, B => position1_N1742, C => n537, D => 
                           n1226, Q => position1_n1490);
   U529 : AOI221 port map( A => n573, B => position1_N2159, C => n571, D => 
                           n1007, Q => position1_n1294);
   U530 : AOI221 port map( A => n540, B => position1_N1744, C => n537, D => 
                           n1224, Q => position1_n1488);
   U531 : AOI221 port map( A => n574, B => position1_N2161, C => n571, D => 
                           n1005, Q => position1_n1292);
   U532 : AOI221 port map( A => n540, B => position1_N1746, C => n537, D => 
                           n1222, Q => position1_n1486);
   U533 : AOI221 port map( A => n574, B => position1_N2163, C => n571, D => 
                           n1003, Q => position1_n1290);
   U534 : AOI221 port map( A => n539, B => position1_N1734, C => n537, D => 
                           n1239, Q => position1_n1498);
   U535 : AOI221 port map( A => n573, B => position1_N2151, C => n571, D => 
                           n1020, Q => position1_n1302);
   U536 : AOI221 port map( A => n539, B => position1_N1736, C => n537, D => 
                           n1235, Q => position1_n1496);
   U537 : AOI221 port map( A => n573, B => position1_N2153, C => n571, D => 
                           n1016, Q => position1_n1300);
   U538 : AOI221 port map( A => n546, B => position1_N1836, C => n545, D => 
                           n1182, Q => position1_n1450);
   U539 : AOI221 port map( A => n580, B => position1_N2253, C => n579, D => 
                           n963, Q => position1_n1254);
   U540 : AOI221 port map( A => n547, B => position1_N1838, C => n545, D => 
                           n1180, Q => position1_n1448);
   U541 : AOI221 port map( A => n581, B => position1_N2255, C => n579, D => 
                           n961, Q => position1_n1252);
   U542 : AOI221 port map( A => n547, B => position1_N1840, C => n545, D => 
                           n1178, Q => position1_n1446);
   U543 : AOI221 port map( A => n581, B => position1_N2257, C => n579, D => 
                           n959, Q => position1_n1250);
   U544 : AOI221 port map( A => n547, B => position1_N1846, C => n545, D => 
                           n1172, Q => position1_n1440);
   U545 : AOI221 port map( A => n581, B => position1_N2263, C => n579, D => 
                           n953, Q => position1_n1244);
   U546 : AOI221 port map( A => n548, B => position1_N1848, C => n545, D => 
                           n1170, Q => position1_n1438);
   U547 : AOI221 port map( A => n582, B => position1_N2265, C => n579, D => 
                           n951, Q => position1_n1242);
   U548 : AOI221 port map( A => n1155, B => n549, C => position1_N1888, D => 
                           n550, Q => position1_n1425);
   U549 : AOI221 port map( A => n936, B => n583, C => position1_N2305, D => 
                           n584, Q => position1_n1229);
   U550 : AOI221 port map( A => n1148, B => n549, C => position1_N1893, D => 
                           n551, Q => position1_n1420);
   U551 : AOI221 port map( A => n929, B => n583, C => position1_N2310, D => 
                           n585, Q => position1_n1224);
   U552 : NOR31 port map( A => position1_N1652, B => position1_N1654, C => 
                           position1_N1653, Q => n1972);
   U553 : NOR31 port map( A => position1_N2069, B => position1_N2071, C => 
                           position1_N2070, Q => n1638);
   U554 : INV3 port map( A => n525, Q => n524);
   U555 : INV3 port map( A => n559, Q => n558);
   U556 : INV3 port map( A => position1_n1521, Q => n1235);
   U557 : AOI221 port map( A => n535, B => position1_N1684, C => n533, D => 
                           position1_N1657, Q => position1_n1521);
   U558 : INV3 port map( A => position1_n1325, Q => n1016);
   U559 : AOI221 port map( A => n569, B => position1_N2101, C => n567, D => 
                           position1_N2074, Q => position1_n1325);
   U560 : INV3 port map( A => position1_n1505, Q => n1216);
   U561 : AOI221 port map( A => n536, B => position1_N1700, C => n533, D => 
                           position1_N1673, Q => position1_n1505);
   U562 : XNR21 port map( A => position1_N1673, B => 
                           position1_sub_216_I4_carry_23_port, Q => 
                           position1_N1700);
   U563 : INV3 port map( A => position1_n1309, Q => n997);
   U564 : AOI221 port map( A => n570, B => position1_N2117, C => n567, D => 
                           position1_N2090, Q => position1_n1309);
   U565 : XNR21 port map( A => position1_N2090, B => 
                           position1_sub_226_I4_carry_23_port, Q => 
                           position1_N2117);
   U566 : NOR21 port map( A => position1_sub_216_I4_carry_23_port, B => 
                           position1_N1673, Q => n116);
   U567 : NOR21 port map( A => position1_sub_226_I4_carry_23_port, B => 
                           position1_N2090, Q => n132);
   U568 : INV3 port map( A => position1_n1449, Q => n1154);
   U569 : AOI221 port map( A => n547, B => position1_N1837, C => n545, D => 
                           n1181, Q => position1_n1449);
   U570 : INV3 port map( A => position1_n1253, Q => n935);
   U571 : AOI221 port map( A => n581, B => position1_N2254, C => n579, D => 
                           n962, Q => position1_n1253);
   U572 : INV3 port map( A => position1_n1518, Q => n1230);
   U573 : AOI221 port map( A => n535, B => position1_N1687, C => n533, D => 
                           position1_N1660, Q => position1_n1518);
   U574 : INV3 port map( A => position1_n1322, Q => n1011);
   U575 : AOI221 port map( A => n569, B => position1_N2104, C => n567, D => 
                           position1_N2077, Q => position1_n1322);
   U576 : INV3 port map( A => position1_n1506, Q => n1217);
   U577 : AOI221 port map( A => n536, B => position1_N1699, C => n533, D => 
                           position1_N1672, Q => position1_n1506);
   U578 : INV3 port map( A => position1_n1310, Q => n998);
   U579 : AOI221 port map( A => n570, B => position1_N2116, C => n567, D => 
                           position1_N2089, Q => position1_n1310);
   U580 : INV3 port map( A => position1_n1484, Q => n1193);
   U581 : AOI221 port map( A => n540, B => position1_N1748, C => n537, D => 
                           n1220, Q => position1_n1484);
   U582 : INV3 port map( A => position1_n1288, Q => n974);
   U583 : AOI221 port map( A => n574, B => position1_N2165, C => n571, D => 
                           n1001, Q => position1_n1288);
   U584 : INV3 port map( A => position1_N1655, Q => n1266);
   U585 : INV3 port map( A => position1_N2072, Q => n1047);
   U586 : INV3 port map( A => position1_n1444, Q => n1146);
   U587 : AOI221 port map( A => n547, B => position1_N1842, C => n545, D => 
                           n1176, Q => position1_n1444);
   U588 : INV3 port map( A => position1_n1248, Q => n927);
   U589 : AOI221 port map( A => n581, B => position1_N2259, C => n579, D => 
                           n957, Q => position1_n1248);
   U590 : INV3 port map( A => position1_n1457, Q => n1164);
   U591 : AOI221 port map( A => n544, B => position1_N1802, C => n541, D => 
                           n1190, Q => position1_n1457);
   U592 : XNR21 port map( A => n1190, B => position1_sub_216_I6_carry_21_port, 
                           Q => position1_N1802);
   U593 : INV3 port map( A => position1_n1261, Q => n945);
   U594 : AOI221 port map( A => n578, B => position1_N2219, C => n575, D => 
                           n971, Q => position1_n1261);
   U595 : XNR21 port map( A => n971, B => position1_sub_226_I6_carry_21_port, Q
                           => position1_N2219);
   U596 : NOR21 port map( A => position1_N1651, B => position1_N1677, Q => 
                           n1973);
   U597 : NOR21 port map( A => position1_N2068, B => position1_N2094, Q => 
                           n1639);
   U598 : INV3 port map( A => position1_n1542, Q => n1290);
   U599 : INV3 port map( A => position1_n1346, Q => n1071);
   U600 : INV3 port map( A => position1_n1540, Q => n1286);
   U601 : INV3 port map( A => position1_n1344, Q => n1067);
   U602 : INV3 port map( A => position1_n1538, Q => n1282);
   U603 : INV3 port map( A => position1_n1342, Q => n1063);
   U604 : INV3 port map( A => position1_n1536, Q => n1278);
   U605 : INV3 port map( A => position1_n1340, Q => n1059);
   U606 : INV3 port map( A => position1_n1534, Q => n1274);
   U607 : INV3 port map( A => position1_n1338, Q => n1055);
   U608 : INV3 port map( A => position1_n1532, Q => n1270);
   U609 : INV3 port map( A => position1_n1336, Q => n1051);
   U610 : INV3 port map( A => position1_n1434, Q => n1132);
   U611 : AOI221 port map( A => n548, B => position1_N1852, C => n545, D => 
                           n1166, Q => position1_n1434);
   U612 : INV3 port map( A => position1_n1238, Q => n913);
   U613 : AOI221 port map( A => n582, B => position1_N2269, C => n579, D => 
                           n947, Q => position1_n1238);
   U614 : INV3 port map( A => position1_n1475, Q => n1182);
   U615 : INV3 port map( A => position1_n1279, Q => n963);
   U616 : INV3 port map( A => position1_n1433, Q => n1131);
   U617 : AOI221 port map( A => n548, B => position1_N1853, C => n545, D => 
                           n1165, Q => position1_n1433);
   U618 : XNR21 port map( A => n1165, B => position1_sub_216_I7_carry_20_port, 
                           Q => position1_N1853);
   U619 : INV3 port map( A => position1_n1237, Q => n912);
   U620 : AOI221 port map( A => n582, B => position1_N2270, C => n579, D => 
                           n946, Q => position1_n1237);
   U621 : XNR21 port map( A => n946, B => position1_sub_226_I7_carry_20_port, Q
                           => position1_N2270);
   U622 : INV3 port map( A => position1_n1481, Q => n1189);
   U623 : AOI221 port map( A => n540, B => position1_N1751, C => n537, D => 
                           n1217, Q => position1_n1481);
   U624 : XNR21 port map( A => n1217, B => position1_sub_216_I5_carry_22_port, 
                           Q => position1_N1751);
   U625 : INV3 port map( A => position1_n1285, Q => n970);
   U626 : AOI221 port map( A => n574, B => position1_N2168, C => n571, D => 
                           n998, Q => position1_n1285);
   U627 : XNR21 port map( A => n998, B => position1_sub_226_I5_carry_22_port, Q
                           => position1_N2168);
   U628 : INV3 port map( A => position1_n1499, Q => n1209);
   U629 : INV3 port map( A => position1_n1303, Q => n990);
   U630 : INV3 port map( A => position1_n1482, Q => n1190);
   U631 : AOI221 port map( A => n540, B => position1_N1750, C => n537, D => 
                           n1218, Q => position1_n1482);
   U632 : INV3 port map( A => position1_n1286, Q => n971);
   U633 : AOI221 port map( A => n574, B => position1_N2167, C => n571, D => 
                           n999, Q => position1_n1286);
   U634 : INV3 port map( A => position1_n1458, Q => n1165);
   U635 : AOI221 port map( A => n544, B => position1_N1801, C => n541, D => 
                           n1191, Q => position1_n1458);
   U636 : INV3 port map( A => position1_n1262, Q => n946);
   U637 : AOI221 port map( A => n578, B => position1_N2218, C => n575, D => 
                           n972, Q => position1_n1262);
   U638 : INV3 port map( A => position1_n1527, Q => n1244);
   U639 : AOI221 port map( A => n534, B => position1_N1651, C => n533, D => 
                           position1_N1651, Q => position1_n1527);
   U640 : INV3 port map( A => position1_n1331, Q => n1025);
   U641 : AOI221 port map( A => n568, B => position1_N2068, C => n567, D => 
                           position1_N2068, Q => position1_n1331);
   U642 : INV3 port map( A => position1_n1528, Q => n1245);
   U643 : AOI221 port map( A => n534, B => position1_N1677, C => n533, D => 
                           position1_N1677, Q => position1_n1528);
   U644 : INV3 port map( A => position1_n1332, Q => n1026);
   U645 : AOI221 port map( A => n568, B => position1_N2094, C => n567, D => 
                           position1_N2094, Q => position1_n1332);
   U646 : INV3 port map( A => position1_n1442, Q => n1144);
   U647 : AOI221 port map( A => n547, B => position1_N1844, C => n545, D => 
                           n1174, Q => position1_n1442);
   U648 : INV3 port map( A => position1_n1246, Q => n925);
   U649 : AOI221 port map( A => n581, B => position1_N2261, C => n579, D => 
                           n955, Q => position1_n1246);
   U650 : INV3 port map( A => position1_n1526, Q => n1243);
   U651 : AOI221 port map( A => n534, B => position1_N1652, C => n533, D => 
                           position1_N1652, Q => position1_n1526);
   U652 : INV3 port map( A => position1_n1330, Q => n1024);
   U653 : AOI221 port map( A => n568, B => position1_N2069, C => n567, D => 
                           position1_N2069, Q => position1_n1330);
   U654 : INV3 port map( A => position1_n1525, Q => n1242);
   U655 : AOI221 port map( A => n534, B => position1_N1653, C => n533, D => 
                           position1_N1653, Q => position1_n1525);
   U656 : INV3 port map( A => position1_n1329, Q => n1023);
   U657 : AOI221 port map( A => n568, B => position1_N2070, C => n567, D => 
                           position1_N2070, Q => position1_n1329);
   U658 : INV3 port map( A => position1_n1504, Q => n1215);
   U659 : AOI221 port map( A => n536, B => position1_N1701, C => n533, D => 
                           position1_N1674, Q => position1_n1504);
   U660 : XNR21 port map( A => position1_sub_216_I4_carry_24_port, B => 
                           position1_N1674, Q => position1_N1701);
   U661 : INV3 port map( A => n116, Q => position1_sub_216_I4_carry_24_port);
   U662 : INV3 port map( A => position1_n1308, Q => n996);
   U663 : AOI221 port map( A => n570, B => position1_N2118, C => n567, D => 
                           position1_N2091, Q => position1_n1308);
   U664 : XNR21 port map( A => position1_sub_226_I4_carry_24_port, B => 
                           position1_N2091, Q => position1_N2118);
   U665 : INV3 port map( A => n132, Q => position1_sub_226_I4_carry_24_port);
   U666 : BUF2 port map( A => position1_N1883, Q => n550);
   U667 : BUF2 port map( A => position1_N2300, Q => n584);
   U668 : INV3 port map( A => position1_n1483, Q => n1191);
   U669 : AOI221 port map( A => n540, B => position1_N1749, C => n537, D => 
                           n1219, Q => position1_n1483);
   U670 : INV3 port map( A => position1_n1287, Q => n972);
   U671 : AOI221 port map( A => n574, B => position1_N2166, C => n571, D => 
                           n1000, Q => position1_n1287);
   U672 : BUF2 port map( A => position1_N1831, Q => n546);
   U673 : BUF2 port map( A => position1_N2248, Q => n580);
   U674 : BUF2 port map( A => position1_N1675, Q => n534);
   U675 : BUF2 port map( A => position1_N2092, Q => n568);
   U676 : BUF2 port map( A => position1_N1727, Q => n538);
   U677 : BUF2 port map( A => position1_N2144, Q => n572);
   U678 : BUF2 port map( A => position1_N1779, Q => n542);
   U679 : BUF2 port map( A => position1_N2196, Q => n576);
   U680 : BUF2 port map( A => position1_N1831, Q => n547);
   U681 : BUF2 port map( A => position1_N2248, Q => n581);
   U682 : BUF2 port map( A => position1_N1675, Q => n535);
   U683 : BUF2 port map( A => position1_N2092, Q => n569);
   U684 : BUF2 port map( A => position1_N1727, Q => n539);
   U685 : BUF2 port map( A => position1_N2144, Q => n573);
   U686 : BUF2 port map( A => position1_N1779, Q => n543);
   U687 : BUF2 port map( A => position1_N2196, Q => n577);
   U688 : BUF2 port map( A => n532, Q => n530);
   U689 : INV3 port map( A => position1_N1623_port, Q => n532);
   U690 : BUF2 port map( A => n566, Q => n564);
   U691 : INV3 port map( A => position1_N2040, Q => n566);
   U692 : BUF2 port map( A => position1_N1883, Q => n551);
   U693 : BUF2 port map( A => position1_N2300, Q => n585);
   U694 : BUF2 port map( A => position1_N1883, Q => n552);
   U695 : BUF2 port map( A => position1_N2300, Q => n586);
   U696 : BUF2 port map( A => position1_N1831, Q => n548);
   U697 : BUF2 port map( A => position1_N2248, Q => n582);
   U698 : BUF2 port map( A => position1_N1675, Q => n536);
   U699 : BUF2 port map( A => position1_N2092, Q => n570);
   U700 : BUF2 port map( A => position1_N1727, Q => n540);
   U701 : BUF2 port map( A => position1_N2144, Q => n574);
   U702 : BUF2 port map( A => position1_N1779, Q => n544);
   U703 : BUF2 port map( A => position1_N2196, Q => n578);
   U704 : INV3 port map( A => n117, Q => position1_sub_216_I5_carry_23_port);
   U705 : NOR21 port map( A => position1_sub_216_I5_carry_22_port, B => n1217, 
                           Q => n117);
   U706 : INV3 port map( A => n133, Q => position1_sub_226_I5_carry_23_port);
   U707 : NOR21 port map( A => position1_sub_226_I5_carry_22_port, B => n998, Q
                           => n133);
   U708 : INV3 port map( A => n119, Q => position1_sub_216_I6_carry_22_port);
   U709 : NOR21 port map( A => position1_sub_216_I6_carry_21_port, B => n1190, 
                           Q => n119);
   U710 : INV3 port map( A => n135, Q => position1_sub_226_I6_carry_22_port);
   U711 : NOR21 port map( A => position1_sub_226_I6_carry_21_port, B => n971, Q
                           => n135);
   U712 : INV3 port map( A => n122, Q => position1_sub_216_I7_carry_21_port);
   U713 : NOR21 port map( A => position1_sub_216_I7_carry_20_port, B => n1165, 
                           Q => n122);
   U714 : INV3 port map( A => n126, Q => position1_sub_216_I8_carry_20_port);
   U715 : NOR21 port map( A => position1_sub_216_I8_carry_19_port, B => n1132, 
                           Q => n126);
   U716 : INV3 port map( A => n138, Q => position1_sub_226_I7_carry_21_port);
   U717 : NOR21 port map( A => position1_sub_226_I7_carry_20_port, B => n946, Q
                           => n138);
   U718 : INV3 port map( A => n142, Q => position1_sub_226_I8_carry_20_port);
   U719 : NOR21 port map( A => position1_sub_226_I8_carry_19_port, B => n913, Q
                           => n142);
   U720 : NOR21 port map( A => n1146, B => n41, Q => n1843);
   U721 : NOR21 port map( A => n927, B => n41, Q => n1509);
   U722 : NAND22 port map( A => n1169, B => n43, Q => n1887);
   U723 : NAND22 port map( A => n950, B => n43, Q => n1553);
   U724 : INV3 port map( A => position1_n1418, Q => n1114);
   U725 : AOI221 port map( A => n1145, B => n549, C => position1_N1895, D => 
                           n551, Q => position1_n1418);
   U726 : INV3 port map( A => position1_n1222, Q => n895);
   U727 : AOI221 port map( A => n926, B => n583, C => position1_N2312, D => 
                           n585, Q => position1_n1222);
   U728 : INV3 port map( A => position1_n1409, Q => n1105);
   U729 : AOI221 port map( A => n1132, B => n549, C => position1_N1904, D => 
                           n552, Q => position1_n1409);
   U730 : XNR21 port map( A => n1132, B => position1_sub_216_I8_carry_19_port, 
                           Q => position1_N1904);
   U731 : INV3 port map( A => position1_n1213, Q => n886);
   U732 : AOI221 port map( A => n913, B => n583, C => position1_N2321, D => 
                           n586, Q => position1_n1213);
   U733 : XNR21 port map( A => n913, B => position1_sub_226_I8_carry_19_port, Q
                           => position1_N2321);
   U734 : INV3 port map( A => position1_n1410, Q => n1106);
   U735 : AOI221 port map( A => n1134, B => n549, C => position1_N1903, D => 
                           n552, Q => position1_n1410);
   U736 : INV3 port map( A => position1_n1214, Q => n887);
   U737 : AOI221 port map( A => n915, B => n583, C => position1_N2320, D => 
                           n586, Q => position1_n1214);
   U738 : BUF2 port map( A => position1_N1883, Q => n553);
   U739 : BUF2 port map( A => position1_N2300, Q => n587);
   U740 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_0_port, Q 
                           => n811);
   U741 : NAND22 port map( A => cam_y_0_port, B => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_0_port);
   U742 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_0_port, Q 
                           => n854);
   U743 : NAND22 port map( A => cam_x_0_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_0_port);
   U744 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_0_port, Q 
                           => n855);
   U745 : NAND22 port map( A => cam_x_0_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_0_port);
   U746 : BUF2 port map( A => n2132, Q => n497);
   U747 : BUF2 port map( A => n2132, Q => cam_x_4_port);
   U748 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_0_port, Q 
                           => n812);
   U749 : NAND22 port map( A => cam_y_0_port, B => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_0_port);
   U750 : BUF2 port map( A => n2130, Q => cam_x_6_port);
   U751 : BUF2 port map( A => n2130, Q => n493);
   U752 : AOI221 port map( A => position1_N606, B => n481, C => position1_N577,
                           D => n480, Q => position1_n1068);
   U753 : XOR21 port map( A => n588, B => position1_r458_carry_17_port, Q => 
                           position1_N577);
   U754 : XOR21 port map( A => position1_r416_carry_17_port, B => n588, Q => 
                           position1_N606);
   U755 : NOR21 port map( A => n300, B => n301, Q => 
                           position1_r458_carry_17_port);
   U756 : INV3 port map( A => position1_n1066, Q => n674);
   U757 : AOI221 port map( A => n635, B => n588, C => position1_n1067, D => 
                           n743, Q => position1_n1066);
   U758 : NAND22 port map( A => position1_n1068, B => position1_n1069, Q => 
                           position1_n1067);
   U759 : AOI221 port map( A => n2, B => n479, C => position1_N447, D => n478, 
                           Q => position1_n1069);
   U760 : XOR21 port map( A => position1_add_250_carry_8_port, B => 
                           position1_dp_cluster_7_N314, Q => position1_N2401);
   U761 : NOR21 port map( A => n313, B => n314, Q => 
                           position1_add_250_carry_8_port);
   U762 : INV3 port map( A => n491, Q => n314);
   U763 : INV3 port map( A => position1_add_250_carry_7_port, Q => n313);
   U764 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, B 
                           => position1_sub_250_3_carry_5_port, Q => 
                           position1_N2387);
   U765 : XNR21 port map( A => n495, B => position1_sub_250_carry_5_port, Q => 
                           position1_N2377);
   U766 : XNR21 port map( A => n491, B => position1_sub_250_carry_7_port, Q => 
                           position1_N2379);
   U767 : NOR21 port map( A => position1_n1056, B => position1_n1057, Q => 
                           position1_n856);
   U768 : XOR21 port map( A => cam_x_2_port, B => 
                           position1_sub_250_carry_2_port, Q => position1_N2374
                           );
   U769 : XOR21 port map( A => n499, B => position1_add_250_carry_3_port, Q => 
                           position1_N2396);
   U770 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, B 
                           => position1_add_250_2_carry_5_port, Q => 
                           position1_N2409);
   U771 : XOR21 port map( A => n495, B => position1_add_250_carry_5_port, Q => 
                           position1_N2398);
   U772 : XOR21 port map( A => n491, B => position1_add_250_carry_7_port, Q => 
                           position1_N2400);
   U773 : NOR40 port map( A => n866, B => position1_n1398, C => cam_x_5_port, D
                           => cam_x_4_port, Q => position1_n1397);
   U774 : INV3 port map( A => position1_n1400, Q => n866);
   U775 : AOI221 port map( A => position1_n1399, B => cam_x_2_port, C => 
                           cam_x_0_port, D => n304, Q => position1_n1398);
   U776 : NOR31 port map( A => cam_x_7_port, B => position1_dp_cluster_7_N314, 
                           C => cam_x_6_port, Q => position1_n1400);
   U777 : XNR21 port map( A => cam_x_3_port, B => 
                           position1_sub_250_carry_3_port, Q => position1_N2375
                           );
   U778 : XNR21 port map( A => n501, B => position1_add_250_carry_2_port, Q => 
                           position1_N2395);
   U779 : NAND41 port map( A => cam_x_5_port, B => cam_x_6_port, C => 
                           cam_x_7_port, D => position1_dp_cluster_7_N314, Q =>
                           position1_n1395);
   U780 : NAND41 port map( A => cam_x_0_port, B => cam_x_1_port, C => n501, D 
                           => cam_x_4_port, Q => position1_n1396);
   U781 : INV3 port map( A => position1_n1397, Q => n853);
   U782 : BUF2 port map( A => position1_n857, Q => n642);
   U783 : BUF2 port map( A => position1_n857, Q => n641);
   U784 : AOI221 port map( A => position1_N537, B => n514, C => 
                           position1_N981_port, D => n642, Q => position1_n946)
                           ;
   U785 : AOI221 port map( A => position1_N538, B => n514, C => 
                           position1_N982_port, D => n642, Q => position1_n942)
                           ;
   U786 : AOI221 port map( A => position1_N539, B => n742, C => 
                           position1_N983_port, D => n642, Q => position1_n938)
                           ;
   U787 : AOI221 port map( A => position1_N540, B => n513, C => 
                           position1_N984_port, D => n642, Q => position1_n934)
                           ;
   U788 : AOI221 port map( A => position1_N487, B => n742, C => 
                           position1_N906_port, D => n643, Q => position1_n1046
                           );
   U789 : AOI221 port map( A => position1_N488, B => n742, C => 
                           position1_N907_port, D => n643, Q => position1_n1042
                           );
   U790 : AOI221 port map( A => position1_N489, B => n742, C => 
                           position1_N908_port, D => n642, Q => position1_n1038
                           );
   U791 : INV3 port map( A => position1_n1179, Q => n714);
   U792 : BUF2 port map( A => position1_n857, Q => n643);
   U793 : INV3 port map( A => position1_n1059, Q => n742);
   U794 : NAND22 port map( A => n743, B => n480, Q => position1_n1059);
   U795 : INV3 port map( A => position1_n1141, Q => n784);
   U796 : INV3 port map( A => n158, Q => position1_add_250_carry_2_port);
   U797 : NOR21 port map( A => cam_x_0_port, B => n503, Q => n158);
   U798 : INV3 port map( A => n148, Q => position1_sub_250_carry_4_port);
   U799 : NOR21 port map( A => position1_sub_250_carry_3_port, B => 
                           cam_x_3_port, Q => n148);
   U800 : INV3 port map( A => n159, Q => position1_add_250_carry_3_port);
   U801 : NOR21 port map( A => position1_add_250_carry_2_port, B => n501, Q => 
                           n159);
   U802 : INV3 port map( A => n155, Q => position1_sub_250_3_carry_6_port);
   U803 : NOR21 port map( A => position1_sub_250_3_carry_5_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, Q 
                           => n155);
   U804 : INV3 port map( A => n150, Q => position1_sub_250_carry_6_port);
   U805 : NOR21 port map( A => position1_sub_250_carry_5_port, B => n495, Q => 
                           n150);
   U806 : INV3 port map( A => position1_N2408, Q => n799);
   U807 : INV3 port map( A => position1_N2410, Q => n791);
   U808 : INV3 port map( A => position1_N2412, Q => n781);
   U809 : INV3 port map( A => position1_N2411, Q => n787);
   U810 : NOR21 port map( A => cam_x_1_port, B => n505, Q => position1_n1399);
   U811 : NOR21 port map( A => n467, B => n302, Q => 
                           position1_sub_250_carry_2_port);
   U812 : INV3 port map( A => n503, Q => n302);
   U813 : NOR21 port map( A => n303, B => n304, Q => 
                           position1_sub_250_carry_3_port);
   U814 : INV3 port map( A => cam_x_2_port, Q => n304);
   U815 : INV3 port map( A => position1_sub_250_carry_2_port, Q => n303);
   U816 : NOR21 port map( A => n309, B => n310, Q => 
                           position1_add_250_carry_6_port);
   U817 : INV3 port map( A => n495, Q => n310);
   U818 : INV3 port map( A => position1_add_250_carry_5_port, Q => n309);
   U819 : NOR21 port map( A => n316, B => gensync1_n94, Q => 
                           position1_add_250_2_carry_6_port);
   U820 : INV3 port map( A => position1_add_250_2_carry_5_port, Q => n316);
   U821 : NOR21 port map( A => n159, B => n306, Q => 
                           position1_add_250_carry_4_port);
   U822 : INV3 port map( A => n499, Q => n306);
   U823 : XOR21 port map( A => n152, B => position1_dp_cluster_7_N314, Q => 
                           position1_N2380);
   U824 : NOR21 port map( A => position1_sub_250_carry_7_port, B => n491, Q => 
                           n152);
   U825 : NOR21 port map( A => position1_n1063, B => position1_n1064, Q => 
                           position1_n859);
   U826 : BUF2 port map( A => n675, Q => n511);
   U827 : BUF2 port map( A => n675, Q => n510);
   U828 : BUF2 port map( A => position1_n858, Q => n645);
   U829 : BUF2 port map( A => position1_n858, Q => n644);
   U830 : BUF2 port map( A => position1_n858, Q => n646);
   U831 : BUF2 port map( A => n675, Q => n512);
   U832 : INV3 port map( A => gensync1_n103, Q => IMG_top_port);
   U833 : INV3 port map( A => position1_r458_carry_16_port, Q => n301);
   U834 : NOR21 port map( A => position1_n1064, B => n484, Q => n482);
   U835 : NOR21 port map( A => position1_n1064, B => n484, Q => n483);
   U836 : NOR21 port map( A => position1_n1064, B => n484, Q => position1_n1154
                           );
   U837 : NAND22 port map( A => image_process1_n57, B => n878, Q => 
                           image_process1_n97);
   U838 : INV3 port map( A => position1_n1064, Q => n743);
   U839 : BUF2 port map( A => position1_n834, Q => n635);
   U840 : INV3 port map( A => position1_n1056, Q => n1361);
   U841 : INV3 port map( A => n589, Q => n588);
   U842 : NAND22 port map( A => image_process1_n113, B => n878, Q => 
                           image_process1_n56);
   U843 : BUF2 port map( A => position1_n834, Q => n636);
   U844 : INV3 port map( A => n2045, Q => n1267);
   U845 : AOI211 port map( A => n2046, B => n2, C => position1_n1530, Q => 
                           n2045);
   U846 : AOI221 port map( A => n2044, B => n2043, C => n45, D => n1269, Q => 
                           n2046);
   U847 : INV3 port map( A => n1711, Q => n1048);
   U848 : AOI211 port map( A => n1712, B => n2, C => position1_n1334, Q => 
                           n1711);
   U849 : AOI221 port map( A => n1710, B => n1709, C => n45, D => n1050, Q => 
                           n1712);
   U850 : INV3 port map( A => position1_N1632_port, Q => n1299);
   U851 : INV3 port map( A => position1_N2049, Q => n1080);
   U852 : XOR21 port map( A => n1301, B => n35, Q => n105);
   U853 : XOR21 port map( A => n1082, B => n35, Q => n106);
   U854 : INV3 port map( A => position1_N1633_port, Q => n1296);
   U855 : INV3 port map( A => position1_N2050, Q => n1077);
   U856 : INV3 port map( A => position1_N1637, Q => n1287);
   U857 : INV3 port map( A => position1_N2054, Q => n1068);
   U858 : INV3 port map( A => position1_N1639, Q => n1283);
   U859 : INV3 port map( A => position1_N2056, Q => n1064);
   U860 : INV3 port map( A => position1_N1641, Q => n1279);
   U861 : INV3 port map( A => position1_N2058, Q => n1060);
   U862 : INV3 port map( A => position1_N1643, Q => n1275);
   U863 : INV3 port map( A => position1_N2060, Q => n1056);
   U864 : INV3 port map( A => position1_N1645, Q => n1271);
   U865 : INV3 port map( A => position1_N2062, Q => n1052);
   U866 : INV3 port map( A => position1_N1635_port, Q => n1291);
   U867 : INV3 port map( A => position1_N2052, Q => n1072);
   U868 : AOI221 port map( A => n526, B => position1_N1582_port, C => n524, D 
                           => position1_N1555_port, Q => position1_n1544);
   U869 : AOI221 port map( A => n560, B => position1_N1999, C => n558, D => 
                           position1_N1972, Q => position1_n1348);
   U870 : XNR21 port map( A => position1_sub_216_I3_carry_24_port, B => 
                           position1_n1529, Q => n107);
   U871 : XNR21 port map( A => position1_sub_226_I3_carry_24_port, B => 
                           position1_n1333, Q => n108);
   U872 : OAI2111 port map( A => n2, B => position1_n1459, C => n1896, D => 
                           n1895, Q => position1_N1831);
   U873 : AOI311 port map( A => n1894, B => n1893, C => n1892, D => n1165, Q =>
                           n1896);
   U874 : NOR40 port map( A => n1161, B => n1162, C => n1163, D => n1164, Q => 
                           n1895);
   U875 : NAND22 port map( A => n588, B => position1_n1459, Q => n1892);
   U876 : OAI2111 port map( A => n2, B => position1_n1263, C => n1562, D => 
                           n1561, Q => position1_N2248);
   U877 : AOI311 port map( A => n1560, B => n1559, C => n1558, D => n946, Q => 
                           n1562);
   U878 : NOR40 port map( A => n942, B => n943, C => n944, D => n945, Q => 
                           n1561);
   U879 : NAND22 port map( A => n588, B => position1_n1263, Q => n1558);
   U880 : OAI2111 port map( A => n2, B => n1246, C => n2009, D => n2008, Q => 
                           position1_N1675);
   U881 : INV3 port map( A => n2007, Q => n1246);
   U882 : NOR21 port map( A => position1_N1674, B => position1_N1673, Q => 
                           n2008);
   U883 : OAI2111 port map( A => n2, B => n1027, C => n1675, D => n1674, Q => 
                           position1_N2092);
   U884 : INV3 port map( A => n1673, Q => n1027);
   U885 : NOR21 port map( A => position1_N2091, B => position1_N2090, Q => 
                           n1674);
   U886 : OAI2111 port map( A => n2, B => n1971, C => n1214, D => n1970, Q => 
                           position1_N1727);
   U887 : INV3 port map( A => n1969, Q => n1214);
   U888 : NOR31 port map( A => n1217, B => n1215, C => n1216, Q => n1970);
   U889 : AOI211 port map( A => n1971, B => n2, C => position1_n1507, Q => 
                           n1969);
   U890 : OAI2111 port map( A => n2, B => n1637, C => n995, D => n1636, Q => 
                           position1_N2144);
   U891 : INV3 port map( A => n1635, Q => n995);
   U892 : NOR31 port map( A => n998, B => n996, C => n997, Q => n1636);
   U893 : AOI211 port map( A => n1637, B => n2, C => position1_n1311, Q => 
                           n1635);
   U894 : OAI2111 port map( A => n2, B => n1934, C => n1933, D => n1932, Q => 
                           position1_N1779);
   U895 : AOI211 port map( A => n1191, B => n1931, C => n1190, Q => n1933);
   U896 : NOR31 port map( A => n1189, B => n1187, C => n1188, Q => n1932);
   U897 : NAND22 port map( A => n588, B => n1934, Q => n1931);
   U898 : OAI2111 port map( A => n2, B => n1600, C => n1599, D => n1598, Q => 
                           position1_N2196);
   U899 : AOI211 port map( A => n972, B => n1597, C => n971, Q => n1599);
   U900 : NOR31 port map( A => n970, B => n968, C => n969, Q => n1598);
   U901 : NAND22 port map( A => n588, B => n1600, Q => n1597);
   U902 : INV3 port map( A => position1_N1647, Q => n1248);
   U903 : INV3 port map( A => position1_N2064, Q => n1029);
   U904 : AOI221 port map( A => n527, B => position1_N1596_port, C => n524, D 
                           => position1_N1569_port, Q => position1_n1530);
   U905 : AOI221 port map( A => n561, B => position1_N2013, C => n558, D => 
                           position1_N1986, Q => position1_n1334);
   U906 : AOI221 port map( A => n526, B => position1_N1584_port, C => n524, D 
                           => position1_N1557_port, Q => position1_n1542);
   U907 : AOI221 port map( A => n560, B => position1_N2001, C => n558, D => 
                           position1_N1974, Q => position1_n1346);
   U908 : AOI221 port map( A => n526, B => position1_N1586_port, C => n524, D 
                           => position1_N1559_port, Q => position1_n1540);
   U909 : AOI221 port map( A => n560, B => position1_N2003, C => n558, D => 
                           position1_N1976, Q => position1_n1344);
   U910 : AOI221 port map( A => n527, B => position1_N1588_port, C => n524, D 
                           => position1_N1561_port, Q => position1_n1538);
   U911 : AOI221 port map( A => n561, B => position1_N2005, C => n558, D => 
                           position1_N1978, Q => position1_n1342);
   U912 : AOI221 port map( A => n527, B => position1_N1590_port, C => n524, D 
                           => position1_N1563_port, Q => position1_n1536);
   U913 : AOI221 port map( A => n561, B => position1_N2007, C => n558, D => 
                           position1_N1980, Q => position1_n1340);
   U914 : AOI221 port map( A => n527, B => position1_N1592_port, C => n524, D 
                           => position1_N1565_port, Q => position1_n1534);
   U915 : AOI221 port map( A => n561, B => position1_N2009, C => n558, D => 
                           position1_N1982, Q => position1_n1338);
   U916 : AOI221 port map( A => n527, B => position1_N1594_port, C => n524, D 
                           => position1_N1567_port, Q => position1_n1532);
   U917 : AOI221 port map( A => n561, B => position1_N2011, C => n558, D => 
                           position1_N1984, Q => position1_n1336);
   U918 : AOI221 port map( A => n539, B => position1_N1733, C => n537, D => 
                           n1241, Q => position1_n1499);
   U919 : XNR21 port map( A => n1241, B => n35, Q => position1_N1733);
   U920 : AOI221 port map( A => n573, B => position1_N2150, C => n571, D => 
                           n1022, Q => position1_n1303);
   U921 : XNR21 port map( A => n1022, B => n35, Q => position1_N2150);
   U922 : AOI221 port map( A => n542, B => position1_N1784, C => n541, D => 
                           n1210, Q => position1_n1475);
   U923 : XNR21 port map( A => n1210, B => n35, Q => position1_N1784);
   U924 : AOI221 port map( A => n576, B => position1_N2201, C => n575, D => 
                           n991, Q => position1_n1279);
   U925 : XNR21 port map( A => n991, B => n35, Q => position1_N2201);
   U926 : NAND22 port map( A => n1859, B => n1858, Q => position1_N1883);
   U927 : NOR40 port map( A => n1131, B => n1132, C => n1857, D => n1856, Q => 
                           n1859);
   U928 : NOR40 port map( A => n1127, B => n1128, C => n1129, D => n1130, Q => 
                           n1858);
   U929 : NOR21 port map( A => n588, B => position1_n1435, Q => n1856);
   U930 : NAND22 port map( A => n1525, B => n1524, Q => position1_N2300);
   U931 : NOR40 port map( A => n912, B => n913, C => n1523, D => n1522, Q => 
                           n1525);
   U932 : NOR40 port map( A => n908, B => n909, C => n910, D => n911, Q => 
                           n1524);
   U933 : NOR21 port map( A => n588, B => position1_n1239, Q => n1522);
   U934 : INV3 port map( A => n523, Q => n522);
   U935 : INV3 port map( A => n557, Q => n556);
   U936 : INV3 port map( A => n523, Q => n521);
   U937 : INV3 port map( A => n557, Q => n555);
   U938 : INV3 port map( A => n523, Q => n520);
   U939 : INV3 port map( A => n557, Q => n554);
   U940 : INV3 port map( A => position1_n1523, Q => n1239);
   U941 : AOI221 port map( A => n535, B => position1_N1682, C => n533, D => 
                           position1_N1655, Q => position1_n1523);
   U942 : XNR21 port map( A => position1_N1655, B => n35, Q => position1_N1682)
                           ;
   U943 : INV3 port map( A => position1_n1327, Q => n1020);
   U944 : AOI221 port map( A => n569, B => position1_N2099, C => n567, D => 
                           position1_N2072, Q => position1_n1327);
   U945 : XNR21 port map( A => position1_N2072, B => n515, Q => position1_N2099
                           );
   U946 : INV3 port map( A => position1_n1451, Q => n1157);
   U947 : AOI221 port map( A => n546, B => position1_N1835, C => n545, D => 
                           n1183, Q => position1_n1451);
   U948 : XNR21 port map( A => n1183, B => n515, Q => position1_N1835);
   U949 : INV3 port map( A => position1_n1255, Q => n938);
   U950 : AOI221 port map( A => n580, B => position1_N2252, C => n579, D => 
                           n964, Q => position1_n1255);
   U951 : XNR21 port map( A => n964, B => n35, Q => position1_N2252);
   U952 : INV3 port map( A => position1_n1547, Q => n1301);
   U953 : INV3 port map( A => position1_n1351, Q => n1082);
   U954 : NAND31 port map( A => position1_n1550, B => position1_n1548, C => 
                           position1_n1549, Q => n109);
   U955 : NAND31 port map( A => position1_n1354, B => position1_n1352, C => 
                           position1_n1353, Q => n110);
   U956 : INV3 port map( A => position1_n1543, Q => n1293);
   U957 : INV3 port map( A => position1_n1347, Q => n1074);
   U958 : INV3 port map( A => position1_n1546, Q => n1300);
   U959 : INV3 port map( A => position1_n1350, Q => n1081);
   U960 : INV3 port map( A => position1_n1541, Q => n1288);
   U961 : INV3 port map( A => position1_n1345, Q => n1069);
   U962 : INV3 port map( A => position1_n1539, Q => n1284);
   U963 : INV3 port map( A => position1_n1343, Q => n1065);
   U964 : INV3 port map( A => position1_n1537, Q => n1280);
   U965 : INV3 port map( A => position1_n1341, Q => n1061);
   U966 : INV3 port map( A => position1_n1535, Q => n1276);
   U967 : INV3 port map( A => position1_n1339, Q => n1057);
   U968 : INV3 port map( A => position1_N1569_port, Q => n1303);
   U969 : INV3 port map( A => position1_N1986, Q => n1084);
   U970 : INV3 port map( A => position1_n1533, Q => n1272);
   U971 : INV3 port map( A => position1_n1337, Q => n1053);
   U972 : INV3 port map( A => position1_n1531, Q => n1269);
   U973 : INV3 port map( A => position1_n1335, Q => n1050);
   U974 : INV3 port map( A => position1_n1334, Q => n1049);
   U975 : INV3 port map( A => position1_n1530, Q => n1268);
   U976 : INV3 port map( A => n168, Q => position1_sub_216_I3_carry_7_port);
   U977 : NOR21 port map( A => n515, B => n1301, Q => n168);
   U978 : INV3 port map( A => n174, Q => position1_sub_226_I3_carry_7_port);
   U979 : NOR21 port map( A => n515, B => n1082, Q => n174);
   U980 : INV3 port map( A => position1_n1545, Q => n1298);
   U981 : INV3 port map( A => position1_n1349, Q => n1079);
   U982 : INV3 port map( A => position1_n1544, Q => n1295);
   U983 : INV3 port map( A => position1_n1348, Q => n1076);
   U984 : INV3 port map( A => n175, Q => position1_sub_226_I4_carry_6_port);
   U985 : NOR21 port map( A => n515, B => position1_N2072, Q => n175);
   U986 : INV3 port map( A => n169, Q => position1_sub_216_I4_carry_6_port);
   U987 : NOR21 port map( A => n515, B => position1_N1655, Q => n169);
   U988 : INV3 port map( A => n170, Q => position1_sub_216_I5_carry_5_port);
   U989 : NOR21 port map( A => n515, B => n1241, Q => n170);
   U990 : INV3 port map( A => n176, Q => position1_sub_226_I5_carry_5_port);
   U991 : NOR21 port map( A => n35, B => n1022, Q => n176);
   U992 : INV3 port map( A => n171, Q => position1_sub_216_I6_carry_4_port);
   U993 : NOR21 port map( A => n515, B => n1210, Q => n171);
   U994 : INV3 port map( A => n177, Q => position1_sub_226_I6_carry_4_port);
   U995 : NOR21 port map( A => n35, B => n991, Q => n177);
   U996 : INV3 port map( A => n172, Q => position1_sub_216_I7_carry_3_port);
   U997 : NOR21 port map( A => n515, B => n1183, Q => n172);
   U998 : INV3 port map( A => n178, Q => position1_sub_226_I7_carry_3_port);
   U999 : NOR21 port map( A => n35, B => n964, Q => n178);
   U1000 : INV3 port map( A => n131, Q => position1_sub_216_I8_carry_2_port);
   U1001 : NOR21 port map( A => n515, B => n1159, Q => n131);
   U1002 : INV3 port map( A => n147, Q => position1_sub_226_I8_carry_2_port);
   U1003 : NOR21 port map( A => n35, B => n940, Q => n147);
   U1004 : NAND31 port map( A => position1_n1553, B => position1_n1551, C => 
                           position1_n1552, Q => n111);
   U1005 : NAND31 port map( A => position1_n1357, B => position1_n1355, C => 
                           position1_n1356, Q => n112);
   U1006 : AOI221 port map( A => n1159, B => n549, C => position1_N1886, D => 
                           n550, Q => position1_n1427);
   U1007 : XNR21 port map( A => n1159, B => n515, Q => position1_N1886);
   U1008 : AOI221 port map( A => n940, B => n583, C => position1_N2303, D => 
                           n584, Q => position1_n1231);
   U1009 : XNR21 port map( A => n940, B => n35, Q => position1_N2303);
   U1010 : BUF2 port map( A => position1_N1571_port, Q => n525);
   U1011 : BUF2 port map( A => position1_N1988, Q => n559);
   U1012 : BUF2 port map( A => position1_N1571_port, Q => n526);
   U1013 : BUF2 port map( A => position1_N1988, Q => n560);
   U1014 : MAJ31 port map( A => position1_n1411, B => n1817, C => n2, Q => 
                           n1821);
   U1015 : AOI221 port map( A => n1107, B => n300, C => n1816, D => n1815, Q =>
                           n1817);
   U1016 : AOI221 port map( A => n1135, B => n549, C => position1_N1902, D => 
                           n552, Q => position1_n1411);
   U1017 : INV3 port map( A => position1_n1412, Q => n1107);
   U1018 : MAJ31 port map( A => position1_n1215, B => n1483, C => n2, Q => 
                           n1487);
   U1019 : AOI221 port map( A => n888, B => n300, C => n1482, D => n1481, Q => 
                           n1483);
   U1020 : AOI221 port map( A => n916, B => n583, C => position1_N2319, D => 
                           n586, Q => position1_n1215);
   U1021 : INV3 port map( A => position1_n1216, Q => n888);
   U1022 : BUF2 port map( A => position1_N1571_port, Q => n527);
   U1023 : BUF2 port map( A => position1_N1988, Q => n561);
   U1024 : NOR21 port map( A => n1157, B => n630, Q => n1828);
   U1025 : NOR21 port map( A => n938, B => n273, Q => n1494);
   U1026 : NOR21 port map( A => n1154, B => n246, Q => n1827);
   U1027 : NOR21 port map( A => n935, B => n246, Q => n1493);
   U1028 : NOR21 port map( A => n1151, B => n278, Q => n1826);
   U1029 : NOR21 port map( A => n932, B => n250, Q => n1492);
   U1030 : NOR21 port map( A => n1142, B => n261, Q => n1825);
   U1031 : NOR21 port map( A => n923, B => n290, Q => n1491);
   U1032 : NOR21 port map( A => n1139, B => n294, Q => n1824);
   U1033 : NOR21 port map( A => n920, B => n265, Q => n1490);
   U1034 : NOR21 port map( A => n1136, B => n269, Q => n1823);
   U1035 : NOR21 port map( A => n917, B => n298, Q => n1489);
   U1036 : NOR21 port map( A => n487, B => n549, Q => position1_N2355);
   U1037 : NOR21 port map( A => n488, B => n583, Q => position1_N2364);
   U1038 : NOR21 port map( A => n489, B => n524, Q => position1_N2361);
   U1039 : NOR21 port map( A => n488, B => n558, Q => position1_N2370);
   U1040 : NOR21 port map( A => n487, B => n533, Q => position1_N2359);
   U1041 : NOR21 port map( A => n487, B => n545, Q => position1_N2356);
   U1042 : NOR21 port map( A => n489, B => n579, Q => position1_N2365);
   U1043 : NOR21 port map( A => n487, B => n537, Q => position1_N2358);
   U1044 : NOR21 port map( A => n487, B => n541, Q => position1_N2357);
   U1045 : NOR21 port map( A => n488, B => n567, Q => position1_N2368);
   U1046 : NOR21 port map( A => n489, B => n571, Q => position1_N2367);
   U1047 : NOR21 port map( A => n488, B => n575, Q => position1_N2366);
   U1048 : INV3 port map( A => n1829, Q => n1158);
   U1049 : AOI211 port map( A => n1160, B => n35, C => n1159, Q => n1829);
   U1050 : INV3 port map( A => n1495, Q => n939);
   U1051 : AOI211 port map( A => n941, B => n35, C => n940, Q => n1495);
   U1052 : NOR21 port map( A => n488, B => n523, Q => position1_N2362);
   U1053 : NOR21 port map( A => n489, B => n557, Q => position1_N2371);
   U1054 : NOR21 port map( A => n489, B => n564, Q => position1_N2369);
   U1055 : NOR21 port map( A => n489, B => n883, Q => position1_N2363);
   U1056 : INV3 port map( A => position1_N2352, Q => n883);
   U1057 : NAND41 port map( A => n1487, B => n1486, C => n1485, D => n1484, Q 
                           => position1_N2352);
   U1058 : NOR21 port map( A => n886, B => n887, Q => n1486);
   U1059 : NOR21 port map( A => n487, B => n530, Q => position1_N2360);
   U1060 : NOR21 port map( A => n487, B => n1102, Q => position1_N2354);
   U1061 : INV3 port map( A => position1_N1935, Q => n1102);
   U1062 : NAND41 port map( A => n1821, B => n1820, C => n1819, D => n1818, Q 
                           => position1_N1935);
   U1063 : NOR21 port map( A => n1105, B => n1106, Q => n1820);
   U1064 : INV3 port map( A => n1936, Q => n1234);
   U1065 : NAND22 port map( A => n274, B => n1235, Q => n1936);
   U1066 : INV3 port map( A => n1602, Q => n1015);
   U1067 : NAND22 port map( A => n274, B => n1016, Q => n1602);
   U1068 : INV3 port map( A => n1938, Q => n1238);
   U1069 : NAND22 port map( A => n630, B => n1239, Q => n1938);
   U1070 : INV3 port map( A => n1604, Q => n1019);
   U1071 : NAND22 port map( A => n630, B => n1020, Q => n1604);
   U1072 : BUF2 port map( A => gensync1_n100, Q => n507);
   U1073 : OAI2111 port map( A => gensync1_N72, B => gensync1_N85, C => n874, D
                           => n871, Q => gensync1_n100);
   U1074 : INV3 port map( A => gensync1_N69, Q => n871);
   U1075 : INV3 port map( A => gensync1_n99, Q => cam_y_0_port);
   U1076 : NOR21 port map( A => n411, B => n412, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_11_port);
   U1077 : INV3 port map( A => position1_N365_port, Q => n412);
   U1078 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_10_port, Q 
                           => n411);
   U1079 : NOR21 port map( A => n349, B => n412, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_11_port);
   U1080 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_10_port, Q 
                           => n349);
   U1081 : NOR21 port map( A => n413, B => n414, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_12_port);
   U1082 : INV3 port map( A => position1_N366_port, Q => n414);
   U1083 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_11_port, Q 
                           => n413);
   U1084 : NOR21 port map( A => n350, B => n414, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_12_port);
   U1085 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_11_port, Q 
                           => n350);
   U1086 : NOR21 port map( A => n439, B => n440, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_12_port);
   U1087 : INV3 port map( A => position1_N291, Q => n440);
   U1088 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_11_port, Q 
                           => n439);
   U1089 : NOR21 port map( A => n366, B => n440, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_12_port);
   U1090 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_11_port, Q 
                           => n366);
   U1091 : NOR21 port map( A => n443, B => n444, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_14_port);
   U1092 : INV3 port map( A => position1_N293, Q => n444);
   U1093 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_13_port, Q 
                           => n443);
   U1094 : NOR21 port map( A => n368, B => n444, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_14_port);
   U1095 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_13_port, Q 
                           => n368);
   U1096 : NOR21 port map( A => n412, B => n231, Q => 
                           position1_r413_carry_11_port);
   U1097 : INV3 port map( A => position1_r413_carry_10_port, Q => n231);
   U1098 : NOR21 port map( A => n416, B => n233, Q => 
                           position1_r413_carry_13_port);
   U1099 : INV3 port map( A => position1_r413_carry_12_port, Q => n233);
   U1100 : NOR21 port map( A => n442, B => n216, Q => 
                           position1_r412_carry_13_port);
   U1101 : INV3 port map( A => position1_r412_carry_12_port, Q => n216);
   U1102 : NOR21 port map( A => n420, B => n235, Q => 
                           position1_r413_carry_15_port);
   U1103 : INV3 port map( A => position1_r413_carry_14_port, Q => n235);
   U1104 : NOR21 port map( A => n446, B => n218, Q => 
                           position1_r412_carry_15_port);
   U1105 : INV3 port map( A => position1_r412_carry_14_port, Q => n218);
   U1106 : NOR21 port map( A => n424, B => n237, Q => 
                           position1_r413_carry_17_port);
   U1107 : INV3 port map( A => position1_r413_carry_16_port, Q => n237);
   U1108 : NOR21 port map( A => n450, B => n220, Q => 
                           position1_r412_carry_17_port);
   U1109 : INV3 port map( A => position1_r412_carry_16_port, Q => n220);
   U1110 : NOR21 port map( A => n428, B => n239, Q => 
                           position1_r413_carry_19_port);
   U1111 : INV3 port map( A => position1_r413_carry_18_port, Q => n239);
   U1112 : NOR21 port map( A => n454, B => n222, Q => 
                           position1_r412_carry_19_port);
   U1113 : INV3 port map( A => position1_r412_carry_18_port, Q => n222);
   U1114 : NOR21 port map( A => n432, B => n241, Q => 
                           position1_r413_carry_21_port);
   U1115 : INV3 port map( A => position1_r413_carry_20_port, Q => n241);
   U1116 : NOR21 port map( A => n458, B => n224, Q => 
                           position1_r412_carry_21_port);
   U1117 : INV3 port map( A => position1_r412_carry_20_port, Q => n224);
   U1118 : NOR21 port map( A => n362, B => n243, Q => 
                           position1_r413_carry_23_port);
   U1119 : INV3 port map( A => position1_r413_carry_22_port, Q => n243);
   U1120 : NOR21 port map( A => n378, B => n226, Q => 
                           position1_r412_carry_23_port);
   U1121 : INV3 port map( A => position1_r412_carry_22_port, Q => n226);
   U1122 : NOR21 port map( A => n414, B => n232, Q => 
                           position1_r413_carry_12_port);
   U1123 : INV3 port map( A => position1_r413_carry_11_port, Q => n232);
   U1124 : NOR21 port map( A => n418, B => n234, Q => 
                           position1_r413_carry_14_port);
   U1125 : INV3 port map( A => position1_r413_carry_13_port, Q => n234);
   U1126 : NOR21 port map( A => n444, B => n217, Q => 
                           position1_r412_carry_14_port);
   U1127 : INV3 port map( A => position1_r412_carry_13_port, Q => n217);
   U1128 : NOR21 port map( A => n422, B => n236, Q => 
                           position1_r413_carry_16_port);
   U1129 : INV3 port map( A => position1_r413_carry_15_port, Q => n236);
   U1130 : NOR21 port map( A => n448, B => n219, Q => 
                           position1_r412_carry_16_port);
   U1131 : INV3 port map( A => position1_r412_carry_15_port, Q => n219);
   U1132 : NOR21 port map( A => n426, B => n238, Q => 
                           position1_r413_carry_18_port);
   U1133 : INV3 port map( A => position1_r413_carry_17_port, Q => n238);
   U1134 : NOR21 port map( A => n452, B => n221, Q => 
                           position1_r412_carry_18_port);
   U1135 : INV3 port map( A => position1_r412_carry_17_port, Q => n221);
   U1136 : NOR21 port map( A => n430, B => n240, Q => 
                           position1_r413_carry_20_port);
   U1137 : INV3 port map( A => position1_r413_carry_19_port, Q => n240);
   U1138 : NOR21 port map( A => n456, B => n223, Q => 
                           position1_r412_carry_20_port);
   U1139 : INV3 port map( A => position1_r412_carry_19_port, Q => n223);
   U1140 : NOR21 port map( A => n434, B => n242, Q => 
                           position1_r413_carry_22_port);
   U1141 : INV3 port map( A => position1_r413_carry_21_port, Q => n242);
   U1142 : NOR21 port map( A => n460, B => n225, Q => 
                           position1_r412_carry_22_port);
   U1143 : INV3 port map( A => position1_r412_carry_21_port, Q => n225);
   U1144 : NOR21 port map( A => n229, B => n230, Q => 
                           position1_r413_carry_10_port);
   U1145 : INV3 port map( A => position1_N364_port, Q => n229);
   U1146 : INV3 port map( A => position1_r413_carry_9_port, Q => n230);
   U1147 : NOR21 port map( A => n212, B => n213, Q => 
                           position1_r412_carry_10_port);
   U1148 : INV3 port map( A => position1_N289, Q => n212);
   U1149 : INV3 port map( A => position1_r412_carry_9_port, Q => n213);
   U1150 : BUF2 port map( A => n2136, Q => n505);
   U1151 : BUF2 port map( A => n2136, Q => cam_x_0_port);
   U1152 : NOR21 port map( A => n228, B => gensync1_n99, Q => 
                           position1_r413_carry_1_port);
   U1153 : INV3 port map( A => position1_N355, Q => n228);
   U1154 : NOR21 port map( A => n211, B => n467, Q => 
                           position1_r412_carry_1_port);
   U1155 : INV3 port map( A => position1_N280, Q => n211);
   U1156 : NOR21 port map( A => n467, B => n466, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_2_port);
   U1157 : INV3 port map( A => position1_N281, Q => n466);
   U1158 : NOR21 port map( A => n467, B => n466, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_2_port);
   U1159 : INV3 port map( A => n505, Q => n467);
   U1160 : NOR21 port map( A => gensync1_n99, B => n468, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_2_port);
   U1161 : INV3 port map( A => position1_N356_port, Q => n468);
   U1162 : NOR21 port map( A => gensync1_n99, B => n468, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_2_port);
   U1163 : XOR21 port map( A => position1_N379, B => 
                           position1_r413_carry_24_port, Q => position1_N559);
   U1164 : NOR21 port map( A => n364, B => n244, Q => 
                           position1_r413_carry_24_port);
   U1165 : INV3 port map( A => position1_r413_carry_23_port, Q => n244);
   U1166 : XOR21 port map( A => position1_N304, B => 
                           position1_r412_carry_24_port, Q => position1_N509);
   U1167 : NOR21 port map( A => n380, B => n227, Q => 
                           position1_r412_carry_24_port);
   U1168 : INV3 port map( A => position1_r412_carry_23_port, Q => n227);
   U1169 : XOR21 port map( A => position1_r412_carry_23_port, B => 
                           position1_N303, Q => position1_N508);
   U1170 : XOR21 port map( A => position1_N303, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_23_port, Q 
                           => position1_N927_port);
   U1171 : BUF2 port map( A => n2135, Q => n503);
   U1172 : BUF2 port map( A => n2135, Q => cam_x_1_port);
   U1173 : NOR21 port map( A => n437, B => n438, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_11_port);
   U1174 : INV3 port map( A => position1_N290, Q => n438);
   U1175 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_10_port, Q 
                           => n437);
   U1176 : NOR21 port map( A => n365, B => n438, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_11_port);
   U1177 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_10_port, Q 
                           => n365);
   U1178 : NOR21 port map( A => n417, B => n418, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_14_port);
   U1179 : INV3 port map( A => position1_N368_port, Q => n418);
   U1180 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_13_port, Q 
                           => n417);
   U1181 : NOR21 port map( A => n352, B => n418, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_14_port);
   U1182 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_13_port, Q 
                           => n352);
   U1183 : NOR21 port map( A => n421, B => n422, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_16_port);
   U1184 : INV3 port map( A => position1_N370_port, Q => n422);
   U1185 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_15_port, Q 
                           => n421);
   U1186 : NOR21 port map( A => n354, B => n422, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_16_port);
   U1187 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_15_port, Q 
                           => n354);
   U1188 : NOR21 port map( A => n447, B => n448, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_16_port);
   U1189 : INV3 port map( A => position1_N295, Q => n448);
   U1190 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_15_port, Q 
                           => n447);
   U1191 : NOR21 port map( A => n370, B => n448, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_16_port);
   U1192 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_15_port, Q 
                           => n370);
   U1193 : NOR21 port map( A => n425, B => n426, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_18_port);
   U1194 : INV3 port map( A => position1_N372, Q => n426);
   U1195 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_17_port, Q 
                           => n425);
   U1196 : NOR21 port map( A => n356, B => n426, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_18_port);
   U1197 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_17_port, Q 
                           => n356);
   U1198 : NOR21 port map( A => n451, B => n452, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_18_port);
   U1199 : INV3 port map( A => position1_N297, Q => n452);
   U1200 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_17_port, Q 
                           => n451);
   U1201 : NOR21 port map( A => n372, B => n452, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_18_port);
   U1202 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_17_port, Q 
                           => n372);
   U1203 : NOR21 port map( A => n429, B => n430, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_20_port);
   U1204 : INV3 port map( A => position1_N374, Q => n430);
   U1205 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_19_port, Q 
                           => n429);
   U1206 : NOR21 port map( A => n358, B => n430, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_20_port);
   U1207 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_19_port, Q 
                           => n358);
   U1208 : NOR21 port map( A => n455, B => n456, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_20_port);
   U1209 : INV3 port map( A => position1_N299, Q => n456);
   U1210 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_19_port, Q 
                           => n455);
   U1211 : NOR21 port map( A => n374, B => n456, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_20_port);
   U1212 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_19_port, Q 
                           => n374);
   U1213 : NOR21 port map( A => n433, B => n434, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_22_port);
   U1214 : INV3 port map( A => position1_N376, Q => n434);
   U1215 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_21_port, Q 
                           => n433);
   U1216 : NOR21 port map( A => n360, B => n434, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_22_port);
   U1217 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_21_port, Q 
                           => n360);
   U1218 : NOR21 port map( A => n459, B => n460, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_22_port);
   U1219 : INV3 port map( A => position1_N301, Q => n460);
   U1220 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_21_port, Q 
                           => n459);
   U1221 : NOR21 port map( A => n376, B => n460, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_22_port);
   U1222 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_21_port, Q 
                           => n376);
   U1223 : NOR21 port map( A => n436, B => n364, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_24_port);
   U1224 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_23_port, Q 
                           => n436);
   U1225 : NOR21 port map( A => n462, B => n380, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_24_port);
   U1226 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_23_port, Q 
                           => n462);
   U1227 : XOR21 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_24_port, B 
                           => position1_N379, Q => position1_N1003_port);
   U1228 : NOR21 port map( A => n363, B => n364, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_24_port);
   U1229 : INV3 port map( A => position1_N378, Q => n364);
   U1230 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_23_port, Q 
                           => n363);
   U1231 : XOR21 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_24_port, B 
                           => position1_N304, Q => position1_N928_port);
   U1232 : NOR21 port map( A => n379, B => n380, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_24_port);
   U1233 : INV3 port map( A => position1_N303, Q => n380);
   U1234 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_23_port, Q 
                           => n379);
   U1235 : NOR21 port map( A => n415, B => n416, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_13_port);
   U1236 : INV3 port map( A => position1_N367_port, Q => n416);
   U1237 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_12_port, Q 
                           => n415);
   U1238 : NOR21 port map( A => n351, B => n416, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_13_port);
   U1239 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_12_port, Q 
                           => n351);
   U1240 : NOR21 port map( A => n441, B => n442, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_13_port);
   U1241 : INV3 port map( A => position1_N292, Q => n442);
   U1242 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_12_port, Q 
                           => n441);
   U1243 : NOR21 port map( A => n367, B => n442, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_13_port);
   U1244 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_12_port, Q 
                           => n367);
   U1245 : NOR21 port map( A => n419, B => n420, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_15_port);
   U1246 : INV3 port map( A => position1_N369_port, Q => n420);
   U1247 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_14_port, Q 
                           => n419);
   U1248 : NOR21 port map( A => n353, B => n420, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_15_port);
   U1249 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_14_port, Q 
                           => n353);
   U1250 : NOR21 port map( A => n445, B => n446, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_15_port);
   U1251 : INV3 port map( A => position1_N294, Q => n446);
   U1252 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_14_port, Q 
                           => n445);
   U1253 : NOR21 port map( A => n369, B => n446, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_15_port);
   U1254 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_14_port, Q 
                           => n369);
   U1255 : NOR21 port map( A => n423, B => n424, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_17_port);
   U1256 : INV3 port map( A => position1_N371, Q => n424);
   U1257 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_16_port, Q 
                           => n423);
   U1258 : NOR21 port map( A => n355, B => n424, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_17_port);
   U1259 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_16_port, Q 
                           => n355);
   U1260 : NOR21 port map( A => n449, B => n450, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_17_port);
   U1261 : INV3 port map( A => position1_N296, Q => n450);
   U1262 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_16_port, Q 
                           => n449);
   U1263 : NOR21 port map( A => n371, B => n450, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_17_port);
   U1264 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_16_port, Q 
                           => n371);
   U1265 : NOR21 port map( A => n427, B => n428, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_19_port);
   U1266 : INV3 port map( A => position1_N373, Q => n428);
   U1267 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_18_port, Q 
                           => n427);
   U1268 : NOR21 port map( A => n357, B => n428, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_19_port);
   U1269 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_18_port, Q 
                           => n357);
   U1270 : NOR21 port map( A => n453, B => n454, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_19_port);
   U1271 : INV3 port map( A => position1_N298, Q => n454);
   U1272 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_18_port, Q 
                           => n453);
   U1273 : NOR21 port map( A => n373, B => n454, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_19_port);
   U1274 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_18_port, Q 
                           => n373);
   U1275 : NOR21 port map( A => n431, B => n432, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_21_port);
   U1276 : INV3 port map( A => position1_N375, Q => n432);
   U1277 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_20_port, Q 
                           => n431);
   U1278 : NOR21 port map( A => n359, B => n432, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_21_port);
   U1279 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_20_port, Q 
                           => n359);
   U1280 : NOR21 port map( A => n457, B => n458, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_21_port);
   U1281 : INV3 port map( A => position1_N300, Q => n458);
   U1282 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_20_port, Q 
                           => n457);
   U1283 : NOR21 port map( A => n375, B => n458, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_21_port);
   U1284 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_20_port, Q 
                           => n375);
   U1285 : NOR21 port map( A => n435, B => n362, Q => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_23_port);
   U1286 : INV3 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_22_port, Q 
                           => n435);
   U1287 : NOR21 port map( A => n361, B => n362, Q => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_23_port);
   U1288 : INV3 port map( A => position1_N377, Q => n362);
   U1289 : INV3 port map( A => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_22_port, Q 
                           => n361);
   U1290 : NOR21 port map( A => n461, B => n378, Q => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_23_port);
   U1291 : INV3 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_22_port, Q 
                           => n461);
   U1292 : NOR21 port map( A => n377, B => n378, Q => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_23_port);
   U1293 : INV3 port map( A => position1_N302, Q => n378);
   U1294 : INV3 port map( A => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_22_port, Q 
                           => n377);
   U1295 : NOR21 port map( A => n440, B => n215, Q => 
                           position1_r412_carry_12_port);
   U1296 : INV3 port map( A => position1_r412_carry_11_port, Q => n215);
   U1297 : NOR21 port map( A => n438, B => n214, Q => 
                           position1_r412_carry_11_port);
   U1298 : INV3 port map( A => position1_r412_carry_10_port, Q => n214);
   U1299 : BUF2 port map( A => n2134, Q => n501);
   U1300 : XOR21 port map( A => position1_r413_carry_23_port, B => 
                           position1_N378, Q => position1_N558);
   U1301 : XOR21 port map( A => position1_r413_carry_22_port, B => 
                           position1_N377, Q => position1_N557);
   U1302 : XOR21 port map( A => position1_r412_carry_21_port, B => 
                           position1_N301, Q => position1_N506);
   U1303 : XOR21 port map( A => position1_r412_carry_22_port, B => 
                           position1_N302, Q => position1_N507);
   U1304 : XOR21 port map( A => position1_N378, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_23_port, Q 
                           => position1_N1002_port);
   U1305 : XOR21 port map( A => position1_N376, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_21_port, Q 
                           => position1_N1000_port);
   U1306 : XOR21 port map( A => position1_N377, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_22_port, Q 
                           => position1_N1001_port);
   U1307 : XOR21 port map( A => position1_N301, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_21_port, Q 
                           => position1_N925_port);
   U1308 : XOR21 port map( A => position1_N302, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_22_port, Q 
                           => position1_N926_port);
   U1309 : BUF2 port map( A => n2134, Q => cam_x_2_port);
   U1310 : BUF2 port map( A => n2133, Q => cam_x_3_port);
   U1311 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_23_port
                           , Q => n410);
   U1312 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_23_port
                           , Q => n395);
   U1313 : INV3 port map( A => position1_n1151, Q => n1363);
   U1314 : INV3 port map( A => position1_n1145, Q => n1362);
   U1315 : XOR21 port map( A => position1_r413_carry_19_port, B => 
                           position1_N374, Q => position1_N554);
   U1316 : XOR21 port map( A => position1_r413_carry_20_port, B => 
                           position1_N375, Q => position1_N555);
   U1317 : XOR21 port map( A => position1_r413_carry_21_port, B => 
                           position1_N376, Q => position1_N556);
   U1318 : XOR21 port map( A => position1_r412_carry_18_port, B => 
                           position1_N298, Q => position1_N503);
   U1319 : XOR21 port map( A => position1_r412_carry_19_port, B => 
                           position1_N299, Q => position1_N504);
   U1320 : XOR21 port map( A => position1_r412_carry_20_port, B => 
                           position1_N300, Q => position1_N505);
   U1321 : XOR21 port map( A => position1_N374, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_19_port, Q 
                           => position1_N998_port);
   U1322 : XOR21 port map( A => position1_N375, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_20_port, Q 
                           => position1_N999_port);
   U1323 : XOR21 port map( A => position1_N298, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_18_port, Q 
                           => position1_N922_port);
   U1324 : XOR21 port map( A => position1_N299, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_19_port, Q 
                           => position1_N923_port);
   U1325 : XOR21 port map( A => position1_N300, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_20_port, Q 
                           => position1_N924_port);
   U1326 : NOR21 port map( A => n507, B => n7, Q => n2132);
   U1327 : BUF2 port map( A => n2133, Q => n499);
   U1328 : INV3 port map( A => gensync1_n94, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port);
   U1329 : NOR21 port map( A => n507, B => n6, Q => n2130);
   U1330 : XOR21 port map( A => position1_r413_carry_17_port, B => 
                           position1_N372, Q => position1_N552);
   U1331 : XOR21 port map( A => position1_r413_carry_18_port, B => 
                           position1_N373, Q => position1_N553);
   U1332 : XOR21 port map( A => position1_r412_carry_16_port, B => 
                           position1_N296, Q => position1_N501);
   U1333 : XOR21 port map( A => position1_r412_carry_17_port, B => 
                           position1_N297, Q => position1_N502);
   U1334 : XOR21 port map( A => position1_N372, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_17_port, Q 
                           => position1_N996_port);
   U1335 : XOR21 port map( A => position1_N373, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_18_port, Q 
                           => position1_N997_port);
   U1336 : XOR21 port map( A => position1_N296, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_16_port, Q 
                           => position1_N920_port);
   U1337 : XOR21 port map( A => position1_N297, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_17_port, Q 
                           => position1_N921_port);
   U1338 : BUF2 port map( A => n2131, Q => n495);
   U1339 : BUF2 port map( A => n2131, Q => cam_x_5_port);
   U1340 : XOR21 port map( A => position1_r413_carry_14_port, B => 
                           position1_N369_port, Q => position1_N549);
   U1341 : XOR21 port map( A => position1_r413_carry_15_port, B => 
                           position1_N370_port, Q => position1_N550);
   U1342 : XOR21 port map( A => position1_r413_carry_16_port, B => 
                           position1_N371, Q => position1_N551);
   U1343 : XOR21 port map( A => position1_r412_carry_14_port, B => 
                           position1_N294, Q => position1_N499);
   U1344 : XOR21 port map( A => position1_r412_carry_15_port, B => 
                           position1_N295, Q => position1_N500);
   U1345 : XOR21 port map( A => position1_N370_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_15_port, Q 
                           => position1_N994_port);
   U1346 : XOR21 port map( A => position1_N371, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_16_port, Q 
                           => position1_N995_port);
   U1347 : XOR21 port map( A => position1_N294, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_14_port, Q 
                           => position1_N918_port);
   U1348 : XOR21 port map( A => position1_N295, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_15_port, Q 
                           => position1_N919_port);
   U1349 : BUF2 port map( A => n2129, Q => cam_x_7_port);
   U1350 : NOR21 port map( A => n507, B => n477, Q => n2128);
   U1351 : XOR21 port map( A => position1_r413_carry_12_port, B => 
                           position1_N367_port, Q => position1_N547);
   U1352 : XOR21 port map( A => position1_r413_carry_13_port, B => 
                           position1_N368_port, Q => position1_N548);
   U1353 : XOR21 port map( A => position1_r412_carry_11_port, B => 
                           position1_N291, Q => position1_N496);
   U1354 : XOR21 port map( A => position1_r412_carry_12_port, B => 
                           position1_N292, Q => position1_N497);
   U1355 : XOR21 port map( A => position1_r412_carry_13_port, B => 
                           position1_N293, Q => position1_N498);
   U1356 : XOR21 port map( A => position1_N367_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_12_port, Q 
                           => position1_N991_port);
   U1357 : XOR21 port map( A => position1_N368_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_13_port, Q 
                           => position1_N992_port);
   U1358 : XOR21 port map( A => position1_N369_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_14_port, Q 
                           => position1_N993_port);
   U1359 : XOR21 port map( A => position1_N292, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_12_port, Q 
                           => position1_N916_port);
   U1360 : XOR21 port map( A => position1_N293, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_13_port, Q 
                           => position1_N917_port);
   U1361 : BUF2 port map( A => n2129, Q => n491);
   U1362 : AOI221 port map( A => position1_N338, B => n646, C => position1_N615
                           , D => n647, Q => position1_n1020);
   U1363 : AOI221 port map( A => position1_N545, B => n514, C => 
                           position1_N989_port, D => n642, Q => position1_n914)
                           ;
   U1364 : XOR21 port map( A => position1_N365_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_10_port, Q 
                           => position1_N989_port);
   U1365 : XOR21 port map( A => position1_r413_carry_10_port, B => 
                           position1_N365_port, Q => position1_N545);
   U1366 : XOR21 port map( A => position1_N365_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_10_port, Q 
                           => position1_N415);
   U1367 : XOR21 port map( A => position1_r413_carry_9_port, B => 
                           position1_N364_port, Q => position1_N544);
   U1368 : XOR21 port map( A => position1_r412_carry_9_port, B => 
                           position1_N289, Q => position1_N494);
   U1369 : XOR21 port map( A => position1_r413_carry_11_port, B => 
                           position1_N366_port, Q => position1_N546);
   U1370 : XOR21 port map( A => position1_r412_carry_10_port, B => 
                           position1_N290, Q => position1_N495);
   U1371 : XOR21 port map( A => position1_N366_port, B => 
                           position1_dp_cluster_2_add_0_root_add_189_3_carry_11_port, Q 
                           => position1_N990_port);
   U1372 : XOR21 port map( A => position1_N290, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_10_port, Q 
                           => position1_N914_port);
   U1373 : XOR21 port map( A => position1_N291, B => 
                           position1_dp_cluster_3_add_0_root_add_188_3_carry_11_port, Q 
                           => position1_N915_port);
   U1374 : INV3 port map( A => position1_n1073, Q => n673);
   U1375 : AOI221 port map( A => n635, B => n595, C => position1_n1074, D => 
                           n743, Q => position1_n1073);
   U1376 : NAND22 port map( A => position1_n1075, B => position1_n1076, Q => 
                           position1_n1074);
   U1377 : AOI221 port map( A => n596, B => n479, C => position1_N446, D => 
                           n478, Q => position1_n1076);
   U1378 : AOI221 port map( A => position1_N412, B => n645, C => position1_N639
                           , D => n649, Q => position1_n924);
   U1379 : AOI221 port map( A => position1_N413, B => n645, C => position1_N640
                           , D => n649, Q => position1_n920);
   U1380 : AOI221 port map( A => position1_N337, B => n646, C => position1_N614
                           , D => n647, Q => position1_n1024);
   U1381 : AOI221 port map( A => position1_N605, B => n481, C => position1_N576
                           , D => n480, Q => position1_n1075);
   U1382 : XOR21 port map( A => position1_r458_carry_16_port, B => n594, Q => 
                           position1_N576);
   U1383 : AOI221 port map( A => position1_N411, B => n645, C => position1_N638
                           , D => n647, Q => position1_n928);
   U1384 : AOI221 port map( A => position1_N335, B => n645, C => position1_N612
                           , D => n647, Q => position1_n1032);
   U1385 : AOI221 port map( A => position1_N336, B => n644, C => position1_N613
                           , D => n647, Q => position1_n1028);
   U1386 : AOI221 port map( A => position1_N603, B => n481, C => position1_N574
                           , D => n480, Q => position1_n1083);
   U1387 : XOR21 port map( A => position1_r458_carry_14_port, B => n476, Q => 
                           position1_N574);
   U1388 : AOI221 port map( A => position1_N604, B => n481, C => position1_N575
                           , D => n480, Q => position1_n1079);
   U1389 : XOR21 port map( A => position1_r458_carry_15_port, B => n598, Q => 
                           position1_N575);
   U1390 : INV3 port map( A => position1_n1081, Q => n671);
   U1391 : AOI221 port map( A => n635, B => position1_N2447, C => 
                           position1_n1082, D => n743, Q => position1_n1081);
   U1392 : NAND22 port map( A => position1_n1083, B => position1_n1084, Q => 
                           position1_n1082);
   U1393 : AOI221 port map( A => position1_N2447, B => n479, C => 
                           position1_N444, D => n478, Q => position1_n1084);
   U1394 : INV3 port map( A => position1_n1077, Q => n672);
   U1395 : AOI221 port map( A => n635, B => n599, C => position1_n1078, D => 
                           n743, Q => position1_n1077);
   U1396 : NAND22 port map( A => position1_n1079, B => position1_n1080, Q => 
                           position1_n1078);
   U1397 : AOI221 port map( A => n600, B => n479, C => position1_N445, D => 
                           n478, Q => position1_n1080);
   U1398 : NAND22 port map( A => reset_top, B => position1_n1182, Q => 
                           position1_n1177);
   U1399 : NAND31 port map( A => position1_n1065, B => position1_n1149, C => 
                           n783, Q => position1_n1063);
   U1400 : INV3 port map( A => position1_n1062, Q => n783);
   U1401 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, B 
                           => position1_add_250_2_carry_4_port, Q => 
                           position1_N2408);
   U1402 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, B 
                           => position1_add_250_2_carry_6_port, Q => 
                           position1_N2410);
   U1403 : XOR21 port map( A => position1_add_250_2_carry_8_port, B => 
                           position1_dp_cluster_6_N389, Q => position1_N2412);
   U1404 : NOR21 port map( A => n318, B => gensync1_n92, Q => 
                           position1_add_250_2_carry_8_port);
   U1405 : INV3 port map( A => position1_add_250_2_carry_7_port, Q => n318);
   U1406 : NAND22 port map( A => position1_n1144, B => position1_n1062, Q => 
                           position1_n1141);
   U1407 : NOR21 port map( A => position1_n1182, B => n653, Q => 
                           position1_n1179);
   U1408 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, B 
                           => position1_sub_250_3_carry_7_port, Q => 
                           position1_N2389);
   U1409 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => position1_add_250_2_carry_3_port, Q => 
                           position1_N2407);
   U1410 : BUF6 port map( A => position1_n1060, Q => n480);
   U1411 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, B 
                           => cam_y_0_port, Q => position1_N2383);
   U1412 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, B 
                           => position1_add_250_2_carry_7_port, Q => 
                           position1_N2411);
   U1413 : NOR21 port map( A => position1_n1057, B => position1_n1058, Q => 
                           position1_n857);
   U1414 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, B 
                           => position1_sub_250_3_carry_4_port, Q => 
                           position1_N2386);
   U1415 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, B 
                           => position1_sub_250_3_carry_6_port, Q => 
                           position1_N2388);
   U1416 : BUF6 port map( A => position1_n1070, Q => n479);
   U1417 : OAI2111 port map( A => n1363, B => position1_n1063, C => 
                           position1_n1142, D => position1_n1143, Q => 
                           position1_n1070);
   U1418 : NAND22 port map( A => position1_n1062, B => n1351, Q => 
                           position1_n1143);
   U1419 : NAND31 port map( A => n784, B => position1_n1145, C => n1361, Q => 
                           position1_n1142);
   U1420 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, B 
                           => position1_add_250_2_carry_2_port, Q => 
                           position1_N2406);
   U1421 : INV3 port map( A => position1_n1085, Q => n670);
   U1422 : AOI221 port map( A => n635, B => n603, C => position1_n1086, D => 
                           n743, Q => position1_n1085);
   U1423 : NAND22 port map( A => position1_n1087, B => position1_n1088, Q => 
                           position1_n1086);
   U1424 : AOI221 port map( A => n604, B => n479, C => position1_N443, D => 
                           n478, Q => position1_n1088);
   U1425 : AOI221 port map( A => n518, B => n479, C => n515, D => n478, Q => 
                           position1_n1140);
   U1426 : AOI221 port map( A => n634, B => n479, C => position1_N431, D => 
                           n478, Q => position1_n1136);
   U1427 : XNR21 port map( A => n517, B => n632, Q => position1_N431);
   U1428 : AOI221 port map( A => n629, B => n479, C => position1_N432, D => 
                           n478, Q => position1_n1132);
   U1429 : XOR21 port map( A => position1_r457_carry_2_port, B => n627, Q => 
                           position1_N432);
   U1430 : AOI221 port map( A => n625, B => n479, C => position1_N433, D => 
                           n478, Q => position1_n1128);
   U1431 : XOR21 port map( A => position1_r457_carry_3_port, B => n623, Q => 
                           position1_N433);
   U1432 : AOI221 port map( A => position1_N2457, B => n479, C => 
                           position1_N434, D => n478, Q => position1_n1124);
   U1433 : XOR21 port map( A => position1_r457_carry_4_port, B => 
                           position1_N2457, Q => position1_N434);
   U1434 : AOI221 port map( A => n622, B => n479, C => position1_N435, D => 
                           n478, Q => position1_n1120);
   U1435 : XOR21 port map( A => position1_r457_carry_5_port, B => n620, Q => 
                           position1_N435);
   U1436 : AOI221 port map( A => n471, B => n479, C => position1_N436, D => 
                           n478, Q => position1_n1116);
   U1437 : XOR21 port map( A => position1_r457_carry_6_port, B => n471, Q => 
                           position1_N436);
   U1438 : AOI221 port map( A => n618, B => n479, C => position1_N437, D => 
                           n478, Q => position1_n1112);
   U1439 : XOR21 port map( A => position1_r457_carry_7_port, B => n615, Q => 
                           position1_N437);
   U1440 : AOI221 port map( A => position1_N2453, B => n479, C => 
                           position1_N438, D => n478, Q => position1_n1108);
   U1441 : XOR21 port map( A => position1_r457_carry_8_port, B => 
                           position1_N2453, Q => position1_N438);
   U1442 : AOI221 port map( A => n612, B => n479, C => position1_N439, D => 
                           n478, Q => position1_n1104);
   U1443 : XOR21 port map( A => position1_r457_carry_9_port, B => n609, Q => 
                           position1_N439);
   U1444 : AOI221 port map( A => n474, B => n479, C => position1_N440, D => 
                           n478, Q => position1_n1100);
   U1445 : XOR21 port map( A => position1_r457_carry_10_port, B => n473, Q => 
                           position1_N440);
   U1446 : AOI221 port map( A => n608, B => n479, C => position1_N441, D => 
                           n478, Q => position1_n1096);
   U1447 : XOR21 port map( A => position1_r457_carry_11_port, B => n606, Q => 
                           position1_N441);
   U1448 : AOI221 port map( A => position1_N2449, B => n479, C => 
                           position1_N442, D => n478, Q => position1_n1092);
   U1449 : XOR21 port map( A => position1_r457_carry_12_port, B => 
                           position1_N2449, Q => position1_N442);
   U1450 : NOR31 port map( A => position1_n1392, B => position1_n1393, C => 
                           position1_n1394, Q => position1_n1391);
   U1451 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, Q 
                           => position1_n1394);
   U1452 : NAND31 port map( A => cam_y_0_port, B => gensync1_n94, C => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, Q 
                           => position1_n1393);
   U1453 : NAND41 port map( A => position1_dp_cluster_6_N389, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, C 
                           => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, D 
                           => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, Q 
                           => position1_n1392);
   U1454 : AOI221 port map( A => position1_N602, B => n481, C => position1_N573
                           , D => n480, Q => position1_n1087);
   U1455 : XOR21 port map( A => position1_r458_carry_13_port, B => n602, Q => 
                           position1_N573);
   U1456 : AOI221 port map( A => position1_N535, B => n513, C => position1_N355
                           , D => n641, Q => position1_n954);
   U1457 : XOR21 port map( A => cam_y_0_port, B => position1_N355, Q => 
                           position1_N535);
   U1458 : AOI221 port map( A => position1_N536, B => n742, C => 
                           position1_N980_port, D => n642, Q => position1_n950)
                           ;
   U1459 : XOR21 port map( A => position1_N356_port, B => cam_y_0_port, Q => 
                           position1_N980_port);
   U1460 : AOI221 port map( A => position1_N485, B => n742, C => position1_N280
                           , D => n641, Q => position1_n1054);
   U1461 : XOR21 port map( A => n505, B => position1_N280, Q => position1_N485)
                           ;
   U1462 : AOI221 port map( A => position1_N486, B => n742, C => 
                           position1_N905_port, D => n643, Q => position1_n1050
                           );
   U1463 : XOR21 port map( A => position1_N281, B => n505, Q => 
                           position1_N905_port);
   U1464 : NOR21 port map( A => position1_N2412, B => n30, Q => n1405);
   U1465 : NOR21 port map( A => position1_N2401, B => n29, Q => n1420);
   U1466 : NOR21 port map( A => position1_N2377, B => n22, Q => n1444);
   U1467 : NOR21 port map( A => position1_N2379, B => n27, Q => n1448);
   U1468 : INV3 port map( A => n153, Q => position1_sub_250_3_carry_4_port);
   U1469 : NOR21 port map( A => position1_sub_250_3_carry_3_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, Q 
                           => n153);
   U1470 : XOR21 port map( A => n157, B => position1_dp_cluster_6_N389, Q => 
                           position1_N2390);
   U1471 : NOR21 port map( A => position1_sub_250_3_carry_7_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, Q 
                           => n157);
   U1472 : INV3 port map( A => n154, Q => position1_sub_250_3_carry_5_port);
   U1473 : NOR21 port map( A => position1_sub_250_3_carry_4_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, Q 
                           => n154);
   U1474 : INV3 port map( A => n160, Q => position1_add_250_2_carry_2_port);
   U1475 : NOR21 port map( A => cam_y_0_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, Q 
                           => n160);
   U1476 : INV3 port map( A => n156, Q => position1_sub_250_3_carry_7_port);
   U1477 : NOR21 port map( A => position1_sub_250_3_carry_6_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, Q 
                           => n156);
   U1478 : INV3 port map( A => position1_n1137, Q => n657);
   U1479 : AOI221 port map( A => n635, B => n517, C => position1_n1138, D => 
                           n743, Q => position1_n1137);
   U1480 : NAND22 port map( A => position1_n1139, B => position1_n1140, Q => 
                           position1_n1138);
   U1481 : AOI221 port map( A => n515, B => n481, C => n519, D => n480, Q => 
                           position1_n1139);
   U1482 : INV3 port map( A => position1_n1133, Q => n658);
   U1483 : AOI221 port map( A => n636, B => n633, C => position1_n1134, D => 
                           n743, Q => position1_n1133);
   U1484 : NAND22 port map( A => position1_n1135, B => position1_n1136, Q => 
                           position1_n1134);
   U1485 : AOI221 port map( A => position1_N590, B => n481, C => n630, D => 
                           n480, Q => position1_n1135);
   U1486 : INV3 port map( A => position1_n1129, Q => n659);
   U1487 : AOI221 port map( A => n636, B => n628, C => position1_n1130, D => 
                           n743, Q => position1_n1129);
   U1488 : NAND22 port map( A => position1_n1131, B => position1_n1132, Q => 
                           position1_n1130);
   U1489 : AOI221 port map( A => position1_N591, B => n481, C => position1_N562
                           , D => n480, Q => position1_n1131);
   U1490 : INV3 port map( A => position1_n1125, Q => n660);
   U1491 : AOI221 port map( A => n636, B => n624, C => position1_n1126, D => 
                           n743, Q => position1_n1125);
   U1492 : NAND22 port map( A => position1_n1127, B => position1_n1128, Q => 
                           position1_n1126);
   U1493 : AOI221 port map( A => position1_N592, B => n481, C => position1_N563
                           , D => n480, Q => position1_n1127);
   U1494 : INV3 port map( A => position1_n1121, Q => n661);
   U1495 : AOI221 port map( A => n636, B => position1_N2457, C => 
                           position1_n1122, D => n743, Q => position1_n1121);
   U1496 : NAND22 port map( A => position1_n1123, B => position1_n1124, Q => 
                           position1_n1122);
   U1497 : AOI221 port map( A => position1_N593, B => n481, C => position1_N564
                           , D => n480, Q => position1_n1123);
   U1498 : INV3 port map( A => position1_n1117, Q => n662);
   U1499 : AOI221 port map( A => n636, B => n621, C => position1_n1118, D => 
                           n743, Q => position1_n1117);
   U1500 : NAND22 port map( A => position1_n1119, B => position1_n1120, Q => 
                           position1_n1118);
   U1501 : AOI221 port map( A => position1_N594, B => n481, C => position1_N565
                           , D => n480, Q => position1_n1119);
   U1502 : INV3 port map( A => position1_n1113, Q => n663);
   U1503 : AOI221 port map( A => n636, B => n471, C => position1_n1114, D => 
                           n743, Q => position1_n1113);
   U1504 : NAND22 port map( A => position1_n1115, B => position1_n1116, Q => 
                           position1_n1114);
   U1505 : AOI221 port map( A => position1_N595, B => n481, C => position1_N566
                           , D => n480, Q => position1_n1115);
   U1506 : INV3 port map( A => position1_n1109, Q => n664);
   U1507 : AOI221 port map( A => n635, B => n617, C => position1_n1110, D => 
                           n743, Q => position1_n1109);
   U1508 : NAND22 port map( A => position1_n1111, B => position1_n1112, Q => 
                           position1_n1110);
   U1509 : AOI221 port map( A => position1_N596, B => n481, C => position1_N567
                           , D => n480, Q => position1_n1111);
   U1510 : INV3 port map( A => position1_n1105, Q => n665);
   U1511 : AOI221 port map( A => n635, B => position1_N2453, C => 
                           position1_n1106, D => n743, Q => position1_n1105);
   U1512 : NAND22 port map( A => position1_n1107, B => position1_n1108, Q => 
                           position1_n1106);
   U1513 : AOI221 port map( A => position1_N597, B => n481, C => position1_N568
                           , D => n480, Q => position1_n1107);
   U1514 : INV3 port map( A => position1_n1101, Q => n666);
   U1515 : AOI221 port map( A => n635, B => n612, C => position1_n1102, D => 
                           n743, Q => position1_n1101);
   U1516 : NAND22 port map( A => position1_n1103, B => position1_n1104, Q => 
                           position1_n1102);
   U1517 : AOI221 port map( A => position1_N598, B => n481, C => position1_N569
                           , D => n480, Q => position1_n1103);
   U1518 : INV3 port map( A => position1_n1097, Q => n667);
   U1519 : AOI221 port map( A => n635, B => n474, C => position1_n1098, D => 
                           n743, Q => position1_n1097);
   U1520 : NAND22 port map( A => position1_n1099, B => position1_n1100, Q => 
                           position1_n1098);
   U1521 : AOI221 port map( A => position1_N599, B => n481, C => position1_N570
                           , D => n480, Q => position1_n1099);
   U1522 : INV3 port map( A => position1_n1093, Q => n668);
   U1523 : AOI221 port map( A => n635, B => n607, C => position1_n1094, D => 
                           n743, Q => position1_n1093);
   U1524 : NAND22 port map( A => position1_n1095, B => position1_n1096, Q => 
                           position1_n1094);
   U1525 : AOI221 port map( A => position1_N600, B => n481, C => position1_N571
                           , D => n480, Q => position1_n1095);
   U1526 : INV3 port map( A => position1_n1089, Q => n669);
   U1527 : AOI221 port map( A => n635, B => position1_N2449, C => 
                           position1_n1090, D => n743, Q => position1_n1089);
   U1528 : NAND22 port map( A => position1_n1091, B => position1_n1092, Q => 
                           position1_n1090);
   U1529 : AOI221 port map( A => position1_N601, B => n481, C => position1_N572
                           , D => n480, Q => position1_n1091);
   U1530 : INV3 port map( A => n161, Q => position1_add_250_2_carry_3_port);
   U1531 : NOR21 port map( A => position1_add_250_2_carry_2_port, B => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, Q 
                           => n161);
   U1532 : NOR21 port map( A => gensync1_n99, B => gensync1_n98, Q => 
                           position1_sub_250_3_carry_2_port);
   U1533 : NOR21 port map( A => n305, B => gensync1_n97, Q => 
                           position1_sub_250_3_carry_3_port);
   U1534 : INV3 port map( A => position1_sub_250_3_carry_2_port, Q => n305);
   U1535 : NOR21 port map( A => n317, B => gensync1_n93, Q => 
                           position1_add_250_2_carry_7_port);
   U1536 : INV3 port map( A => position1_add_250_2_carry_6_port, Q => n317);
   U1537 : NOR21 port map( A => n315, B => gensync1_n95, Q => 
                           position1_add_250_2_carry_5_port);
   U1538 : INV3 port map( A => position1_add_250_2_carry_4_port, Q => n315);
   U1539 : NOR21 port map( A => n161, B => gensync1_n96, Q => 
                           position1_add_250_2_carry_4_port);
   U1540 : NOR31 port map( A => position1_n1064, B => position1_n1062, C => 
                           position1_n1065, Q => position1_n858);
   U1541 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, B 
                           => position1_sub_250_3_carry_2_port, Q => 
                           position1_N2384);
   U1542 : BUF6 port map( A => position1_n1072, Q => n481);
   U1543 : INV3 port map( A => position1_n1061, Q => n675);
   U1544 : AOI311 port map( A => n743, B => n1351, C => position1_n1062, D => 
                           n635, Q => position1_n1061);
   U1545 : NOR21 port map( A => n250, B => n251, Q => 
                           position1_r457_carry_6_port);
   U1546 : INV3 port map( A => n620, Q => n250);
   U1547 : INV3 port map( A => position1_r457_carry_5_port, Q => n251);
   U1548 : NOR21 port map( A => n256, B => n257, Q => 
                           position1_r457_carry_9_port);
   U1549 : INV3 port map( A => position1_N2453, Q => n256);
   U1550 : INV3 port map( A => position1_r457_carry_8_port, Q => n257);
   U1551 : NOR21 port map( A => n286, B => n258, Q => 
                           position1_r457_carry_10_port);
   U1552 : INV3 port map( A => position1_r457_carry_9_port, Q => n258);
   U1553 : NOR21 port map( A => n269, B => n270, Q => 
                           position1_r457_carry_16_port);
   U1554 : INV3 port map( A => n598, Q => n269);
   U1555 : INV3 port map( A => position1_r457_carry_15_port, Q => n270);
   U1556 : NOR21 port map( A => n248, B => n249, Q => 
                           position1_r457_carry_5_port);
   U1557 : INV3 port map( A => position1_N2457, Q => n248);
   U1558 : INV3 port map( A => position1_r457_carry_4_port, Q => n249);
   U1559 : NOR21 port map( A => n246, B => n247, Q => 
                           position1_r457_carry_4_port);
   U1560 : INV3 port map( A => n623, Q => n246);
   U1561 : INV3 port map( A => position1_r457_carry_3_port, Q => n247);
   U1562 : NOR21 port map( A => n245, B => n115, Q => 
                           position1_r457_carry_3_port);
   U1563 : INV3 port map( A => n627, Q => n245);
   U1564 : XOR21 port map( A => n588, B => position1_r457_carry_17_port, Q => 
                           position1_N447);
   U1565 : NOR21 port map( A => n300, B => n271, Q => 
                           position1_r457_carry_17_port);
   U1566 : INV3 port map( A => position1_r457_carry_16_port, Q => n271);
   U1567 : XOR21 port map( A => position1_r457_carry_16_port, B => n594, Q => 
                           position1_N446);
   U1568 : INV3 port map( A => n115, Q => position1_r457_carry_2_port);
   U1569 : NOR21 port map( A => n632, B => n517, Q => n115);
   U1570 : NOR21 port map( A => n265, B => n266, Q => 
                           position1_r457_carry_14_port);
   U1571 : INV3 port map( A => n602, Q => n265);
   U1572 : INV3 port map( A => position1_r457_carry_13_port, Q => n266);
   U1573 : NOR21 port map( A => n261, B => n262, Q => 
                           position1_r457_carry_12_port);
   U1574 : INV3 port map( A => n606, Q => n261);
   U1575 : INV3 port map( A => position1_r457_carry_11_port, Q => n262);
   U1576 : NOR21 port map( A => n252, B => n253, Q => 
                           position1_r457_carry_7_port);
   U1577 : INV3 port map( A => n471, Q => n252);
   U1578 : INV3 port map( A => position1_r457_carry_6_port, Q => n253);
   U1579 : NOR21 port map( A => n263, B => n264, Q => 
                           position1_r457_carry_13_port);
   U1580 : INV3 port map( A => n475, Q => n263);
   U1581 : INV3 port map( A => position1_r457_carry_12_port, Q => n264);
   U1582 : NOR21 port map( A => n267, B => n268, Q => 
                           position1_r457_carry_15_port);
   U1583 : INV3 port map( A => position1_N2447, Q => n267);
   U1584 : INV3 port map( A => position1_r457_carry_14_port, Q => n268);
   U1585 : NOR21 port map( A => n254, B => n255, Q => 
                           position1_r457_carry_8_port);
   U1586 : INV3 port map( A => n615, Q => n254);
   U1587 : INV3 port map( A => position1_r457_carry_7_port, Q => n255);
   U1588 : NOR21 port map( A => n259, B => n260, Q => 
                           position1_r457_carry_11_port);
   U1589 : INV3 port map( A => n473, Q => n259);
   U1590 : INV3 port map( A => position1_r457_carry_10_port, Q => n260);
   U1591 : NAND41 port map( A => n874, B => gensync1_n104, C => n816, D => 
                           gensync1_N85, Q => gensync1_n103);
   U1592 : NOR21 port map( A => gensync1_N69, B => gensync1_N72, Q => 
                           gensync1_n104);
   U1593 : NOR21 port map( A => n272, B => n273, Q => 
                           position1_r458_carry_3_port);
   U1594 : INV3 port map( A => n632, Q => n273);
   U1595 : INV3 port map( A => n627, Q => n272);
   U1596 : NOR21 port map( A => n274, B => n275, Q => 
                           position1_r458_carry_4_port);
   U1597 : INV3 port map( A => n623, Q => n274);
   U1598 : INV3 port map( A => position1_r458_carry_3_port, Q => n275);
   U1599 : NOR21 port map( A => n276, B => n277, Q => 
                           position1_r458_carry_5_port);
   U1600 : INV3 port map( A => n469, Q => n276);
   U1601 : INV3 port map( A => position1_r458_carry_4_port, Q => n277);
   U1602 : NOR21 port map( A => n280, B => n281, Q => 
                           position1_r458_carry_7_port);
   U1603 : INV3 port map( A => n470, Q => n280);
   U1604 : INV3 port map( A => position1_r458_carry_6_port, Q => n281);
   U1605 : NOR21 port map( A => n286, B => n287, Q => 
                           position1_r458_carry_10_port);
   U1606 : INV3 port map( A => n609, Q => n286);
   U1607 : INV3 port map( A => position1_r458_carry_9_port, Q => n287);
   U1608 : NOR21 port map( A => n288, B => n289, Q => 
                           position1_r458_carry_11_port);
   U1609 : INV3 port map( A => n473, Q => n288);
   U1610 : INV3 port map( A => position1_r458_carry_10_port, Q => n289);
   U1611 : XOR21 port map( A => position1_N356_port, B => cam_y_0_port, Q => 
                           position1_N406);
   U1612 : XOR21 port map( A => position1_N281, B => n505, Q => position1_N331)
                           ;
   U1613 : XOR21 port map( A => position1_r457_carry_14_port, B => 
                           position1_N2447, Q => position1_N444);
   U1614 : XOR21 port map( A => position1_r457_carry_15_port, B => n598, Q => 
                           position1_N445);
   U1615 : NOR21 port map( A => n294, B => n295, Q => 
                           position1_r458_carry_14_port);
   U1616 : INV3 port map( A => n602, Q => n294);
   U1617 : INV3 port map( A => position1_r458_carry_13_port, Q => n295);
   U1618 : NOR21 port map( A => n298, B => n299, Q => 
                           position1_r458_carry_16_port);
   U1619 : INV3 port map( A => n598, Q => n298);
   U1620 : INV3 port map( A => position1_r458_carry_15_port, Q => n299);
   U1621 : NOR21 port map( A => n278, B => n279, Q => 
                           position1_r458_carry_6_port);
   U1622 : INV3 port map( A => n620, Q => n278);
   U1623 : INV3 port map( A => position1_r458_carry_5_port, Q => n279);
   U1624 : NOR21 port map( A => n290, B => n291, Q => 
                           position1_r458_carry_12_port);
   U1625 : INV3 port map( A => n606, Q => n290);
   U1626 : INV3 port map( A => position1_r458_carry_11_port, Q => n291);
   U1627 : NOR21 port map( A => n282, B => n283, Q => 
                           position1_r458_carry_8_port);
   U1628 : INV3 port map( A => n615, Q => n282);
   U1629 : INV3 port map( A => position1_r458_carry_7_port, Q => n283);
   U1630 : NOR21 port map( A => n292, B => n293, Q => 
                           position1_r458_carry_13_port);
   U1631 : INV3 port map( A => n475, Q => n292);
   U1632 : INV3 port map( A => position1_r458_carry_12_port, Q => n293);
   U1633 : NOR21 port map( A => n296, B => n297, Q => 
                           position1_r458_carry_15_port);
   U1634 : INV3 port map( A => n476, Q => n296);
   U1635 : INV3 port map( A => position1_r458_carry_14_port, Q => n297);
   U1636 : NOR21 port map( A => n284, B => n285, Q => 
                           position1_r458_carry_9_port);
   U1637 : INV3 port map( A => n472, Q => n284);
   U1638 : INV3 port map( A => position1_r458_carry_8_port, Q => n285);
   U1639 : NOR21 port map( A => image_process1_n117, B => gensync1_n103, Q => 
                           image_process1_n57);
   U1640 : XOR21 port map( A => position1_r457_carry_13_port, B => n602, Q => 
                           position1_N443);
   U1641 : NOR41 port map( A => n777, B => image_process1_N59_port, C => 
                           image_process1_N62_port, D => 
                           image_process1_N64_port, Q => image_process1_n89);
   U1642 : INV3 port map( A => image_process1_n57, Q => n777);
   U1643 : NOR21 port map( A => gensync1_n103, B => n776, Q => 
                           image_process1_n58);
   U1644 : INV3 port map( A => image_process1_n117, Q => n776);
   U1645 : NAND22 port map( A => gensync1_n103, B => position1_n1176, Q => 
                           position1_n1175);
   U1646 : NOR21 port map( A => image_process1_n97, B => 
                           image_process1_N62_port, Q => image_process1_n95);
   U1647 : XOR21 port map( A => position1_r458_carry_11_port, B => n606, Q => 
                           position1_N571);
   U1648 : XOR21 port map( A => position1_r458_carry_12_port, B => n475, Q => 
                           position1_N572);
   U1649 : INV3 port map( A => n490, Q => n815);
   U1650 : BUF2 port map( A => n484, Q => n485);
   U1651 : AOI211 port map( A => n489, B => position1_n1175, C => n655, Q => 
                           n484);
   U1652 : NOR21 port map( A => n509, B => n820, Q => gensync1_N63);
   U1653 : INV3 port map( A => gensync1_N53, Q => n820);
   U1654 : NOR21 port map( A => n509, B => n819, Q => gensync1_N64);
   U1655 : INV3 port map( A => gensync1_N54, Q => n819);
   U1656 : NOR21 port map( A => gensync1_n102, B => n828, Q => gensync1_N30);
   U1657 : INV3 port map( A => gensync1_N20, Q => n828);
   U1658 : XOR21 port map( A => position1_r458_carry_8_port, B => n472, Q => 
                           position1_N568);
   U1659 : XOR21 port map( A => position1_r458_carry_9_port, B => n609, Q => 
                           position1_N569);
   U1660 : XOR21 port map( A => position1_r458_carry_10_port, B => n473, Q => 
                           position1_N570);
   U1661 : INV3 port map( A => position1_n1144, Q => n1351);
   U1662 : NOR21 port map( A => gensync1_n102, B => n829, Q => gensync1_N29);
   U1663 : INV3 port map( A => gensync1_N19, Q => n829);
   U1664 : NOR21 port map( A => gensync1_n102, B => n830, Q => gensync1_N28);
   U1665 : INV3 port map( A => gensync1_N18, Q => n830);
   U1666 : NOR21 port map( A => n509, B => n821, Q => gensync1_N62);
   U1667 : INV3 port map( A => gensync1_N52, Q => n821);
   U1668 : NOR21 port map( A => n509, B => n822, Q => gensync1_N61);
   U1669 : INV3 port map( A => gensync1_N51, Q => n822);
   U1670 : NAND22 port map( A => position1_n1176, B => n650, Q => 
                           position1_n1064);
   U1671 : INV3 port map( A => n656, Q => n650);
   U1672 : NAND22 port map( A => position1_n1058, B => position1_n1146, Q => 
                           position1_n1056);
   U1673 : NOR21 port map( A => n652, B => n488, Q => position1_n834);
   U1674 : XOR21 port map( A => position1_r458_carry_6_port, B => n470, Q => 
                           position1_N566);
   U1675 : XOR21 port map( A => position1_r458_carry_7_port, B => n615, Q => 
                           position1_N567);
   U1676 : NOR21 port map( A => gensync1_n102, B => n831, Q => gensync1_N27);
   U1677 : INV3 port map( A => gensync1_N17, Q => n831);
   U1678 : BUF2 port map( A => position1_n1152, Q => n488);
   U1679 : NOR21 port map( A => n508, B => n823, Q => gensync1_N60);
   U1680 : INV3 port map( A => gensync1_N50, Q => n823);
   U1681 : NOR21 port map( A => image_process1_n113, B => 
                           image_process1_N59_port, Q => image_process1_n112);
   U1682 : INV3 port map( A => image_process1_N59_port, Q => n878);
   U1683 : XOR21 port map( A => position1_r458_carry_3_port, B => n623, Q => 
                           position1_N563);
   U1684 : XOR21 port map( A => position1_r458_carry_4_port, B => n469, Q => 
                           position1_N564);
   U1685 : XOR21 port map( A => position1_r458_carry_5_port, B => n620, Q => 
                           position1_N565);
   U1686 : BUF2 port map( A => position1_n1152, Q => n489);
   U1687 : NOR21 port map( A => gensync1_n102, B => n832, Q => gensync1_N26);
   U1688 : INV3 port map( A => gensync1_N16, Q => n832);
   U1689 : NOR21 port map( A => gensync1_n102, B => n833, Q => gensync1_N25);
   U1690 : INV3 port map( A => gensync1_N15, Q => n833);
   U1691 : BUF2 port map( A => n102, Q => n589);
   U1692 : NOR21 port map( A => n877, B => image_process1_N62_port, Q => 
                           image_process1_n113);
   U1693 : INV3 port map( A => image_process1_N64_port, Q => n877);
   U1694 : BUF2 port map( A => gensync1_n101, Q => n509);
   U1695 : BUF2 port map( A => gensync1_n101, Q => n508);
   U1696 : INV3 port map( A => gensync1_N129, Q => n817);
   U1697 : NOR21 port map( A => n508, B => n824, Q => gensync1_N59);
   U1698 : INV3 port map( A => gensync1_N49, Q => n824);
   U1699 : NOR21 port map( A => n508, B => n825, Q => gensync1_N58);
   U1700 : INV3 port map( A => gensync1_N48, Q => n825);
   U1701 : NOR21 port map( A => n508, B => n826, Q => gensync1_N57);
   U1702 : INV3 port map( A => gensync1_N47, Q => n826);
   U1703 : INV3 port map( A => n654, Q => n651);
   U1704 : XOR21 port map( A => n632, B => n627, Q => position1_N562);
   U1705 : NOR21 port map( A => gensync1_n102, B => n834, Q => gensync1_N24);
   U1706 : INV3 port map( A => gensync1_N14, Q => n834);
   U1707 : NOR21 port map( A => gensync1_n102, B => n835, Q => gensync1_N23);
   U1708 : INV3 port map( A => gensync1_N13, Q => n835);
   U1709 : INV3 port map( A => n631, Q => n630);
   U1710 : INV3 port map( A => n516, Q => n515);
   U1711 : INV3 port map( A => n594, Q => n300);
   U1712 : INV3 port map( A => position1_N1570_port, Q => n1302);
   U1713 : AOI221 port map( A => position1_N1569_port, B => n45, C => n2081, D 
                           => n2080, Q => n2082);
   U1714 : NAND22 port map( A => n595, B => n1303, Q => n2080);
   U1715 : INV3 port map( A => position1_N1987, Q => n1083);
   U1716 : AOI221 port map( A => position1_N1986, B => n300, C => n1747, D => 
                           n1746, Q => n1748);
   U1717 : NAND22 port map( A => n595, B => n1084, Q => n1746);
   U1718 : NAND22 port map( A => position1_N1530_port, B => n521, Q => 
                           position1_n1569);
   U1719 : NAND22 port map( A => position1_N1947, B => n555, Q => 
                           position1_n1373);
   U1720 : NAND22 port map( A => position1_N1532_port, B => n521, Q => 
                           position1_n1567);
   U1721 : NAND22 port map( A => position1_N1949, B => n555, Q => 
                           position1_n1371);
   U1722 : NAND22 port map( A => position1_N1534_port, B => n520, Q => 
                           position1_n1565);
   U1723 : NAND22 port map( A => position1_N1951, B => n554, Q => 
                           position1_n1369);
   U1724 : NAND22 port map( A => position1_N1536_port, B => n520, Q => 
                           position1_n1563);
   U1725 : NAND22 port map( A => position1_N1953, B => n554, Q => 
                           position1_n1367);
   U1726 : NAND22 port map( A => position1_N1538_port, B => n520, Q => 
                           position1_n1561);
   U1727 : NAND22 port map( A => position1_N1955, B => n554, Q => 
                           position1_n1365);
   U1728 : NAND22 port map( A => position1_N1540_port, B => n520, Q => 
                           position1_n1559);
   U1729 : NAND22 port map( A => position1_N1957, B => n554, Q => 
                           position1_n1363);
   U1730 : NAND22 port map( A => position1_N1542_port, B => n520, Q => 
                           position1_n1557);
   U1731 : NAND22 port map( A => position1_N1959, B => n554, Q => 
                           position1_n1361);
   U1732 : NAND22 port map( A => position1_N1544_port, B => n520, Q => 
                           position1_n1555);
   U1733 : NAND22 port map( A => position1_N1961, B => n554, Q => 
                           position1_n1359);
   U1734 : AOI221 port map( A => n526, B => position1_N1581_port, C => n524, D 
                           => position1_N1554_port, Q => position1_n1545);
   U1735 : AOI221 port map( A => n560, B => position1_N1998, C => n558, D => 
                           position1_N1971, Q => position1_n1349);
   U1736 : AOI221 port map( A => n526, B => position1_N1580_port, C => n524, D 
                           => position1_N1553_port, Q => position1_n1546);
   U1737 : XNR21 port map( A => position1_N1553_port, B => n515, Q => 
                           position1_N1580_port);
   U1738 : AOI221 port map( A => n560, B => position1_N1997, C => n558, D => 
                           position1_N1970, Q => position1_n1350);
   U1739 : XNR21 port map( A => position1_N1970, B => n515, Q => 
                           position1_N1997);
   U1740 : AOI221 port map( A => n526, B => position1_N1585_port, C => n524, D 
                           => position1_N1558_port, Q => position1_n1541);
   U1741 : AOI221 port map( A => n560, B => position1_N2002, C => n558, D => 
                           position1_N1975, Q => position1_n1345);
   U1742 : AOI221 port map( A => n526, B => position1_N1587_port, C => n524, D 
                           => position1_N1560_port, Q => position1_n1539);
   U1743 : AOI221 port map( A => n560, B => position1_N2004, C => n558, D => 
                           position1_N1977, Q => position1_n1343);
   U1744 : AOI221 port map( A => n527, B => position1_N1589_port, C => n524, D 
                           => position1_N1562_port, Q => position1_n1537);
   U1745 : AOI221 port map( A => n561, B => position1_N2006, C => n558, D => 
                           position1_N1979, Q => position1_n1341);
   U1746 : AOI221 port map( A => n527, B => position1_N1591_port, C => n524, D 
                           => position1_N1564_port, Q => position1_n1535);
   U1747 : AOI221 port map( A => n561, B => position1_N2008, C => n558, D => 
                           position1_N1981, Q => position1_n1339);
   U1748 : AOI221 port map( A => n527, B => position1_N1593_port, C => n524, D 
                           => position1_N1566_port, Q => position1_n1533);
   U1749 : AOI221 port map( A => n561, B => position1_N2010, C => n558, D => 
                           position1_N1983, Q => position1_n1337);
   U1750 : AOI221 port map( A => n527, B => position1_N1595_port, C => n524, D 
                           => position1_N1568_port, Q => position1_n1531);
   U1751 : AOI221 port map( A => n561, B => position1_N2012, C => n558, D => 
                           position1_N1985, Q => position1_n1335);
   U1752 : AOI221 port map( A => n527, B => position1_N1597_port, C => n524, D 
                           => position1_N1570_port, Q => position1_n1529);
   U1753 : AOI221 port map( A => n561, B => position1_N2014, C => n558, D => 
                           position1_N1987, Q => position1_n1333);
   U1754 : AOI221 port map( A => n526, B => position1_N1552_port, C => n524, D 
                           => position1_N1552_port, Q => position1_n1547);
   U1755 : AOI221 port map( A => n560, B => position1_N1969, C => n558, D => 
                           position1_N1969, Q => position1_n1351);
   U1756 : AOI221 port map( A => n526, B => position1_N1550_port, C => n524, D 
                           => position1_N1550_port, Q => position1_n1549);
   U1757 : AOI221 port map( A => n525, B => position1_N1549_port, C => n524, D 
                           => position1_N1549_port, Q => position1_n1550);
   U1758 : AOI221 port map( A => n560, B => position1_N1967, C => n558, D => 
                           position1_N1967, Q => position1_n1353);
   U1759 : AOI221 port map( A => n559, B => position1_N1966, C => n558, D => 
                           position1_N1966, Q => position1_n1354);
   U1760 : AOI221 port map( A => n526, B => position1_N1551_port, C => n524, D 
                           => position1_N1551_port, Q => position1_n1548);
   U1761 : AOI221 port map( A => n560, B => position1_N1968, C => n558, D => 
                           position1_N1968, Q => position1_n1352);
   U1762 : AOI221 port map( A => n525, B => position1_N1547_port, C => n524, D 
                           => position1_N1547_port, Q => position1_n1552);
   U1763 : AOI221 port map( A => n525, B => position1_N1548_port, C => n524, D 
                           => position1_N1548_port, Q => position1_n1551);
   U1764 : AOI221 port map( A => n525, B => position1_N1573_port, C => n524, D 
                           => position1_N1573_port, Q => position1_n1553);
   U1765 : AOI221 port map( A => n559, B => position1_N1964, C => n558, D => 
                           position1_N1964, Q => position1_n1356);
   U1766 : AOI221 port map( A => n559, B => position1_N1965, C => n558, D => 
                           position1_N1965, Q => position1_n1355);
   U1767 : AOI221 port map( A => n559, B => position1_N1990, C => n558, D => 
                           position1_N1990, Q => position1_n1357);
   U1768 : INV3 port map( A => position1_N1671, Q => n1249);
   U1769 : NOR21 port map( A => position1_N1671, B => n45, Q => n2006);
   U1770 : INV3 port map( A => position1_N2088, Q => n1030);
   U1771 : NOR21 port map( A => position1_N2088, B => n300, Q => n1672);
   U1772 : AOI221 port map( A => n526, B => position1_N1583_port, C => n524, D 
                           => position1_N1556_port, Q => position1_n1543);
   U1773 : AOI221 port map( A => n560, B => position1_N2000, C => n558, D => 
                           position1_N1973, Q => position1_n1347);
   U1774 : AOI221 port map( A => n1192, B => n1930, C => n45, D => n1193, Q => 
                           n1934);
   U1775 : INV3 port map( A => n1897, Q => n1192);
   U1776 : AOI221 port map( A => position1_n1485, B => n599, C => n1186, D => 
                           n1195, Q => n1930);
   U1777 : NOR21 port map( A => n1193, B => n300, Q => n1897);
   U1778 : AOI221 port map( A => n973, B => n1596, C => n45, D => n974, Q => 
                           n1600);
   U1779 : INV3 port map( A => n1563, Q => n973);
   U1780 : AOI221 port map( A => position1_n1289, B => n599, C => n967, D => 
                           n976, Q => n1596);
   U1781 : NOR21 port map( A => n974, B => n300, Q => n1563);
   U1782 : OAI2111 port map( A => position1_n1436, B => n596, C => n1854, D => 
                           n1853, Q => n1855);
   U1783 : NAND22 port map( A => n298, B => n1136, Q => n1854);
   U1784 : OAI2111 port map( A => n296, B => n1137, C => n1126, D => n1852, Q 
                           => n1853);
   U1785 : INV3 port map( A => n1823, Q => n1126);
   U1786 : OAI2111 port map( A => position1_n1240, B => n596, C => n1520, D => 
                           n1519, Q => n1521);
   U1787 : NAND22 port map( A => n269, B => n917, Q => n1520);
   U1788 : OAI2111 port map( A => n267, B => n918, C => n907, D => n1518, Q => 
                           n1519);
   U1789 : INV3 port map( A => n1489, Q => n907);
   U1790 : OAI2111 port map( A => position1_n1254, B => n629, C => n1497, D => 
                           n1496, Q => n1498);
   U1791 : NAND22 port map( A => n273, B => n938, Q => n1497);
   U1792 : OAI2111 port map( A => n35, B => n941, C => n937, D => n939, Q => 
                           n1496);
   U1793 : INV3 port map( A => n1494, Q => n937);
   U1794 : OAI2111 port map( A => position1_n1252, B => position1_N2457, C => 
                           n1500, D => n1499, Q => n1501);
   U1795 : NAND22 port map( A => n246, B => n935, Q => n1500);
   U1796 : OAI2111 port map( A => n67, B => n936, C => n934, D => n1498, Q => 
                           n1499);
   U1797 : INV3 port map( A => n1493, Q => n934);
   U1798 : OAI2111 port map( A => position1_n1250, B => n471, C => n1503, D => 
                           n1502, Q => n1504);
   U1799 : NAND22 port map( A => n278, B => n932, Q => n1503);
   U1800 : OAI2111 port map( A => n248, B => n933, C => n931, D => n1501, Q => 
                           n1502);
   U1801 : INV3 port map( A => n1492, Q => n931);
   U1802 : OAI2111 port map( A => position1_n1440, B => n475, C => n1848, D => 
                           n1847, Q => n1849);
   U1803 : NAND22 port map( A => n261, B => n1142, Q => n1848);
   U1804 : OAI2111 port map( A => n259, B => n1144, C => n1141, D => n1143, Q 
                           => n1847);
   U1805 : INV3 port map( A => n1825, Q => n1141);
   U1806 : OAI2111 port map( A => position1_n1244, B => position1_N2449, C => 
                           n1514, D => n1513, Q => n1515);
   U1807 : NAND22 port map( A => n290, B => n923, Q => n1514);
   U1808 : OAI2111 port map( A => n259, B => n925, C => n922, D => n924, Q => 
                           n1513);
   U1809 : INV3 port map( A => n1491, Q => n922);
   U1810 : OAI2111 port map( A => position1_n1446, B => n470, C => n1837, D => 
                           n1836, Q => n1838);
   U1811 : NAND22 port map( A => n250, B => n1151, Q => n1837);
   U1812 : OAI2111 port map( A => n276, B => n1152, C => n1150, D => n1835, Q 
                           => n1836);
   U1813 : INV3 port map( A => n1826, Q => n1150);
   U1814 : OAI2111 port map( A => position1_n1438, B => n476, C => n1851, D => 
                           n1850, Q => n1852);
   U1815 : NAND22 port map( A => n294, B => n1139, Q => n1851);
   U1816 : OAI2111 port map( A => n292, B => n1140, C => n1138, D => n1849, Q 
                           => n1850);
   U1817 : INV3 port map( A => n1824, Q => n1138);
   U1818 : OAI2111 port map( A => position1_n1242, B => position1_N2447, C => 
                           n1517, D => n1516, Q => n1518);
   U1819 : NAND22 port map( A => n265, B => n920, Q => n1517);
   U1820 : OAI2111 port map( A => n263, B => n921, C => n919, D => n1515, Q => 
                           n1516);
   U1821 : INV3 port map( A => n1490, Q => n919);
   U1822 : OAI2111 port map( A => position1_n1448, B => n469, C => n1834, D => 
                           n1833, Q => n1835);
   U1823 : NAND22 port map( A => n274, B => n1154, Q => n1834);
   U1824 : OAI2111 port map( A => n67, B => n1155, C => n1153, D => n1832, Q =>
                           n1833);
   U1825 : INV3 port map( A => n1827, Q => n1153);
   U1826 : OAI2111 port map( A => position1_n1450, B => n629, C => n1831, D => 
                           n1830, Q => n1832);
   U1827 : NAND22 port map( A => n273, B => n1157, Q => n1831);
   U1828 : OAI2111 port map( A => n515, B => n1160, C => n1156, D => n1158, Q 
                           => n1830);
   U1829 : INV3 port map( A => n1828, Q => n1156);
   U1830 : INV3 port map( A => n1939, Q => n1240);
   U1831 : NOR40 port map( A => n1242, B => n1243, C => n1244, D => n1245, Q =>
                           n1940);
   U1832 : NAND22 port map( A => position1_n1524, B => n517, Q => n1939);
   U1833 : INV3 port map( A => n1605, Q => n1021);
   U1834 : NOR40 port map( A => n1023, B => n1024, C => n1025, D => n1026, Q =>
                           n1606);
   U1835 : NAND22 port map( A => position1_n1328, B => n517, Q => n1605);
   U1836 : NOR21 port map( A => n624, B => position1_n1544, Q => n2018);
   U1837 : INV3 port map( A => n2010, Q => n1297);
   U1838 : NOR21 port map( A => n623, B => position1_n1348, Q => n1684);
   U1839 : INV3 port map( A => n1676, Q => n1078);
   U1840 : INV3 port map( A => n1937, Q => n1236);
   U1841 : NAND22 port map( A => position1_n1522, B => n627, Q => n1937);
   U1842 : INV3 port map( A => n1603, Q => n1017);
   U1843 : NAND22 port map( A => position1_n1326, B => n627, Q => n1603);
   U1844 : INV3 port map( A => n1935, Q => n1232);
   U1845 : NAND22 port map( A => position1_n1520, B => n469, Q => n1935);
   U1846 : INV3 port map( A => n1601, Q => n1013);
   U1847 : NAND22 port map( A => position1_n1324, B => position1_N2457, Q => 
                           n1601);
   U1848 : AOI2111 port map( A => n595, B => position1_n1436, C => n1133, D => 
                           n1125, Q => n1857);
   U1849 : INV3 port map( A => n1822, Q => n1133);
   U1850 : INV3 port map( A => n1855, Q => n1125);
   U1851 : NAND22 port map( A => position1_n1435, B => n588, Q => n1822);
   U1852 : AOI2111 port map( A => n593, B => position1_n1240, C => n914, D => 
                           n906, Q => n1523);
   U1853 : INV3 port map( A => n1488, Q => n914);
   U1854 : INV3 port map( A => n1521, Q => n906);
   U1855 : NAND22 port map( A => position1_n1239, B => n588, Q => n1488);
   U1856 : AOI221 port map( A => n1968, B => n1967, C => n45, D => n1219, Q => 
                           n1971);
   U1857 : NAND22 port map( A => position1_n1508, B => n594, Q => n1968);
   U1858 : AOI221 port map( A => position1_n1509, B => n599, C => n1966, D => 
                           n1965, Q => n1967);
   U1859 : NAND22 port map( A => n68, B => n1220, Q => n1966);
   U1860 : AOI221 port map( A => n1634, B => n1633, C => n45, D => n1000, Q => 
                           n1637);
   U1861 : NAND22 port map( A => position1_n1312, B => n594, Q => n1634);
   U1862 : AOI221 port map( A => position1_n1313, B => n597, C => n1632, D => 
                           n1631, Q => n1633);
   U1863 : NAND22 port map( A => n298, B => n1001, Q => n1632);
   U1864 : NOR21 port map( A => n1210, B => n35, Q => n1899);
   U1865 : NOR31 port map( A => n1213, B => n1211, C => n1212, Q => n1900);
   U1866 : NOR21 port map( A => n991, B => n35, Q => n1565);
   U1867 : NOR31 port map( A => n994, B => n992, C => n993, Q => n1566);
   U1868 : NOR21 port map( A => n1208, B => n272, Q => n1904);
   U1869 : NOR21 port map( A => n632, B => position1_n1499, Q => n1902);
   U1870 : NOR21 port map( A => n989, B => n245, Q => n1570);
   U1871 : NOR21 port map( A => n632, B => position1_n1303, Q => n1568);
   U1872 : NOR21 port map( A => n1206, B => n276, Q => n1908);
   U1873 : NOR21 port map( A => n623, B => position1_n1497, Q => n1906);
   U1874 : NOR21 port map( A => n987, B => n42, Q => n1574);
   U1875 : NOR21 port map( A => n623, B => position1_n1301, Q => n1572);
   U1876 : NOR21 port map( A => n1204, B => n46, Q => n1912);
   U1877 : NOR21 port map( A => n621, B => position1_n1495, Q => n1910);
   U1878 : NOR21 port map( A => n985, B => n252, Q => n1578);
   U1879 : NOR21 port map( A => n620, B => position1_n1299, Q => n1576);
   U1880 : NOR21 port map( A => n1202, B => n284, Q => n1916);
   U1881 : NOR21 port map( A => n616, B => position1_n1493, Q => n1914);
   U1882 : NOR21 port map( A => n983, B => n41, Q => n1582);
   U1883 : NOR21 port map( A => n615, B => position1_n1297, Q => n1580);
   U1884 : NOR21 port map( A => n1200, B => n47, Q => n1920);
   U1885 : NOR21 port map( A => n610, B => position1_n1491, Q => n1918);
   U1886 : NOR21 port map( A => n981, B => n288, Q => n1586);
   U1887 : NOR21 port map( A => n610, B => position1_n1295, Q => n1584);
   U1888 : AOI221 port map( A => position1_n1542, B => n622, C => n2022, D => 
                           n2021, Q => n2023);
   U1889 : NAND22 port map( A => n278, B => n1290, Q => n2022);
   U1890 : AOI221 port map( A => n2020, B => n1292, C => n248, D => n1293, Q =>
                           n2021);
   U1891 : INV3 port map( A => n2019, Q => n1292);
   U1892 : AOI221 port map( A => position1_n1346, B => n619, C => n1688, D => 
                           n1687, Q => n1689);
   U1893 : NAND22 port map( A => n250, B => n1071, Q => n1688);
   U1894 : AOI221 port map( A => n1686, B => n1073, C => n248, D => n1074, Q =>
                           n1687);
   U1895 : INV3 port map( A => n1685, Q => n1073);
   U1896 : AOI221 port map( A => position1_n1540, B => n617, C => n2026, D => 
                           n2025, Q => n2027);
   U1897 : NAND22 port map( A => n282, B => n1286, Q => n2026);
   U1898 : AOI221 port map( A => n2024, B => n2023, C => n280, D => n1288, Q =>
                           n2025);
   U1899 : NAND22 port map( A => position1_n1541, B => n470, Q => n2024);
   U1900 : AOI221 port map( A => position1_n1344, B => n617, C => n1692, D => 
                           n1691, Q => n1693);
   U1901 : NAND22 port map( A => n254, B => n1067, Q => n1692);
   U1902 : AOI221 port map( A => n1690, B => n1689, C => n252, D => n1069, Q =>
                           n1691);
   U1903 : NAND22 port map( A => position1_n1345, B => n471, Q => n1690);
   U1904 : AOI221 port map( A => position1_n1538, B => n612, C => n2030, D => 
                           n2029, Q => n2031);
   U1905 : NAND22 port map( A => n286, B => n1282, Q => n2030);
   U1906 : AOI221 port map( A => n2028, B => n2027, C => n284, D => n1284, Q =>
                           n2029);
   U1907 : NAND22 port map( A => position1_n1539, B => n472, Q => n2028);
   U1908 : AOI221 port map( A => position1_n1342, B => n611, C => n1696, D => 
                           n1695, Q => n1697);
   U1909 : NAND22 port map( A => n286, B => n1063, Q => n1696);
   U1910 : AOI221 port map( A => n1694, B => n1693, C => n256, D => n1065, Q =>
                           n1695);
   U1911 : NAND22 port map( A => position1_n1343, B => n472, Q => n1694);
   U1912 : AOI221 port map( A => position1_n1536, B => n607, C => n2034, D => 
                           n2033, Q => n2035);
   U1913 : NAND22 port map( A => n39, B => n1278, Q => n2034);
   U1914 : AOI221 port map( A => n2032, B => n2031, C => n288, D => n1280, Q =>
                           n2033);
   U1915 : NAND22 port map( A => position1_n1537, B => n473, Q => n2032);
   U1916 : AOI221 port map( A => position1_n1340, B => n605, C => n1700, D => 
                           n1699, Q => n1701);
   U1917 : NAND22 port map( A => n261, B => n1059, Q => n1700);
   U1918 : AOI221 port map( A => n1698, B => n1697, C => n288, D => n1061, Q =>
                           n1699);
   U1919 : NAND22 port map( A => position1_n1341, B => n473, Q => n1698);
   U1920 : NOR21 port map( A => n1198, B => n44, Q => n1924);
   U1921 : NOR21 port map( A => n606, B => position1_n1489, Q => n1922);
   U1922 : NOR21 port map( A => n979, B => n263, Q => n1590);
   U1923 : NOR21 port map( A => n606, B => position1_n1293, Q => n1588);
   U1924 : AOI221 port map( A => position1_n1534, B => n603, C => n2038, D => 
                           n2037, Q => n2039);
   U1925 : NAND22 port map( A => n40, B => n1274, Q => n2038);
   U1926 : AOI221 port map( A => n2036, B => n2035, C => n292, D => n1276, Q =>
                           n2037);
   U1927 : NAND22 port map( A => position1_n1535, B => n475, Q => n2036);
   U1928 : AOI221 port map( A => position1_n1338, B => n601, C => n1704, D => 
                           n1703, Q => n1705);
   U1929 : NAND22 port map( A => n294, B => n1055, Q => n1704);
   U1930 : AOI221 port map( A => n1702, B => n1701, C => n292, D => n1057, Q =>
                           n1703);
   U1931 : NAND22 port map( A => position1_n1339, B => n475, Q => n1702);
   U1932 : AOI221 port map( A => position1_n1532, B => n599, C => n2042, D => 
                           n2041, Q => n2043);
   U1933 : NAND22 port map( A => n68, B => n1270, Q => n2042);
   U1934 : AOI221 port map( A => n2040, B => n2039, C => n267, D => n1272, Q =>
                           n2041);
   U1935 : NAND22 port map( A => position1_n1533, B => n476, Q => n2040);
   U1936 : AOI221 port map( A => position1_n1336, B => n599, C => n1708, D => 
                           n1707, Q => n1709);
   U1937 : NAND22 port map( A => n269, B => n1051, Q => n1708);
   U1938 : AOI221 port map( A => n1706, B => n1705, C => n296, D => n1053, Q =>
                           n1707);
   U1939 : NAND22 port map( A => position1_n1337, B => n476, Q => n1706);
   U1940 : INV3 port map( A => position1_N1659, Q => n1262);
   U1941 : NOR21 port map( A => position1_N1659, B => n248, Q => n1982);
   U1942 : INV3 port map( A => position1_N2076, Q => n1043);
   U1943 : NOR21 port map( A => position1_N2076, B => n42, Q => n1648);
   U1944 : INV3 port map( A => position1_N1657, Q => n1264);
   U1945 : NOR21 port map( A => position1_N1657, B => n272, Q => n1978);
   U1946 : INV3 port map( A => position1_N2074, Q => n1045);
   U1947 : NOR21 port map( A => position1_N2074, B => n245, Q => n1644);
   U1948 : INV3 port map( A => position1_N1661, Q => n1260);
   U1949 : NOR21 port map( A => position1_N1661, B => n46, Q => n1986);
   U1950 : INV3 port map( A => position1_N2078, Q => n1041);
   U1951 : NOR21 port map( A => position1_N2078, B => n252, Q => n1652);
   U1952 : INV3 port map( A => position1_N1663, Q => n1258);
   U1953 : NOR21 port map( A => position1_N1663, B => n256, Q => n1990);
   U1954 : INV3 port map( A => position1_N2080, Q => n1039);
   U1955 : NOR21 port map( A => position1_N2080, B => n41, Q => n1656);
   U1956 : INV3 port map( A => position1_N1665, Q => n1256);
   U1957 : NOR21 port map( A => position1_N1665, B => n47, Q => n1994);
   U1958 : INV3 port map( A => position1_N2082, Q => n1037);
   U1959 : NOR21 port map( A => position1_N2082, B => n288, Q => n1660);
   U1960 : INV3 port map( A => position1_N1667, Q => n1254);
   U1961 : NOR21 port map( A => position1_N1667, B => n44, Q => n1998);
   U1962 : INV3 port map( A => position1_N2084, Q => n1035);
   U1963 : NOR21 port map( A => position1_N2084, B => n292, Q => n1664);
   U1964 : INV3 port map( A => position1_N1669, Q => n1252);
   U1965 : NOR21 port map( A => position1_N1669, B => n43, Q => n2002);
   U1966 : INV3 port map( A => position1_N2086, Q => n1033);
   U1967 : NOR21 port map( A => position1_N2086, B => n296, Q => n1668);
   U1968 : AOI221 port map( A => n2048, B => n2047, C => n518, D => n1304, Q =>
                           n2049);
   U1969 : INV3 port map( A => position1_N1553_port, Q => n1304);
   U1970 : NOR31 port map( A => position1_N1573_port, B => position1_N1548_port
                           , C => position1_N1547_port, Q => n2048);
   U1971 : NOR40 port map( A => position1_N1552_port, B => position1_N1551_port
                           , C => position1_N1550_port, D => 
                           position1_N1549_port, Q => n2047);
   U1972 : AOI221 port map( A => n1714, B => n1713, C => n518, D => n1085, Q =>
                           n1715);
   U1973 : INV3 port map( A => position1_N1970, Q => n1085);
   U1974 : NOR31 port map( A => position1_N1990, B => position1_N1965, C => 
                           position1_N1964, Q => n1714);
   U1975 : NOR40 port map( A => position1_N1969, B => position1_N1968, C => 
                           position1_N1967, D => position1_N1966, Q => n1713);
   U1976 : AOI221 port map( A => n1168, B => n269, C => n1890, D => n1889, Q =>
                           n1891);
   U1977 : NAND22 port map( A => n600, B => position1_n1461, Q => n1889);
   U1978 : AOI221 port map( A => n1888, B => n1887, C => n476, D => 
                           position1_n1462, Q => n1890);
   U1979 : AOI221 port map( A => n949, B => n298, C => n1556, D => n1555, Q => 
                           n1557);
   U1980 : NAND22 port map( A => n600, B => position1_n1265, Q => n1555);
   U1981 : AOI221 port map( A => n1554, B => n1553, C => position1_N2447, D => 
                           position1_n1266, Q => n1556);
   U1982 : AOI2111 port map( A => n1146, B => n256, C => n1841, D => n1147, Q 
                           => n1842);
   U1983 : INV3 port map( A => n1840, Q => n1147);
   U1984 : NOR21 port map( A => n616, B => position1_n1445, Q => n1841);
   U1985 : OAI2111 port map( A => n280, B => n1149, C => n1839, D => n1838, Q 
                           => n1840);
   U1986 : AOI2111 port map( A => n927, B => n284, C => n1507, D => n928, Q => 
                           n1508);
   U1987 : INV3 port map( A => n1506, Q => n928);
   U1988 : NOR21 port map( A => n615, B => position1_n1249, Q => n1507);
   U1989 : OAI2111 port map( A => n252, B => n930, C => n1505, D => n1504, Q =>
                           n1506);
   U1990 : AOI221 port map( A => n1952, B => n1951, C => n284, D => n1227, Q =>
                           n1953);
   U1991 : NAND22 port map( A => position1_n1516, B => position1_N2453, Q => 
                           n1952);
   U1992 : AOI221 port map( A => position1_n1517, B => n617, C => n1950, D => 
                           n1949, Q => n1951);
   U1993 : NAND22 port map( A => n282, B => n1228, Q => n1950);
   U1994 : AOI221 port map( A => n1618, B => n1617, C => n256, D => n1008, Q =>
                           n1619);
   U1995 : NAND22 port map( A => position1_n1320, B => position1_N2453, Q => 
                           n1618);
   U1996 : AOI221 port map( A => position1_n1321, B => n615, C => n1616, D => 
                           n1615, Q => n1617);
   U1997 : NAND22 port map( A => n254, B => n1009, Q => n1616);
   U1998 : AOI221 port map( A => n1956, B => n1955, C => n259, D => n1225, Q =>
                           n1957);
   U1999 : NAND22 port map( A => position1_n1514, B => n473, Q => n1956);
   U2000 : AOI221 port map( A => position1_n1515, B => n612, C => n1954, D => 
                           n1953, Q => n1955);
   U2001 : NAND22 port map( A => n286, B => n1226, Q => n1954);
   U2002 : AOI221 port map( A => n1622, B => n1621, C => n288, D => n1006, Q =>
                           n1623);
   U2003 : NAND22 port map( A => position1_n1318, B => n473, Q => n1622);
   U2004 : AOI221 port map( A => position1_n1319, B => n611, C => n1620, D => 
                           n1619, Q => n1621);
   U2005 : NAND22 port map( A => n286, B => n1007, Q => n1620);
   U2006 : AOI221 port map( A => n1960, B => n1959, C => n263, D => n1223, Q =>
                           n1961);
   U2007 : NAND22 port map( A => position1_n1512, B => position1_N2449, Q => 
                           n1960);
   U2008 : AOI221 port map( A => position1_n1513, B => n607, C => n1958, D => 
                           n1957, Q => n1959);
   U2009 : NAND22 port map( A => n39, B => n1224, Q => n1958);
   U2010 : AOI221 port map( A => n1626, B => n1625, C => n292, D => n1004, Q =>
                           n1627);
   U2011 : NAND22 port map( A => position1_n1316, B => position1_N2449, Q => 
                           n1626);
   U2012 : AOI221 port map( A => position1_n1317, B => n607, C => n1624, D => 
                           n1623, Q => n1625);
   U2013 : NAND22 port map( A => n290, B => n1005, Q => n1624);
   U2014 : AOI221 port map( A => n1964, B => n1963, C => n267, D => n1221, Q =>
                           n1965);
   U2015 : NAND22 port map( A => position1_n1510, B => position1_N2447, Q => 
                           n1964);
   U2016 : AOI221 port map( A => position1_n1511, B => n603, C => n1962, D => 
                           n1961, Q => n1963);
   U2017 : NAND22 port map( A => n40, B => n1222, Q => n1962);
   U2018 : AOI221 port map( A => n1630, B => n1629, C => n296, D => n1002, Q =>
                           n1631);
   U2019 : NAND22 port map( A => position1_n1314, B => position1_N2447, Q => 
                           n1630);
   U2020 : AOI221 port map( A => position1_n1315, B => n603, C => n1628, D => 
                           n1627, Q => n1629);
   U2021 : NAND22 port map( A => n265, B => n1003, Q => n1628);
   U2022 : AOI221 port map( A => n1948, B => n1229, C => n280, D => n1230, Q =>
                           n1949);
   U2023 : INV3 port map( A => n1947, Q => n1229);
   U2024 : NAND22 port map( A => position1_n1519, B => n621, Q => n1948);
   U2025 : AOI221 port map( A => n1614, B => n1010, C => n252, D => n1011, Q =>
                           n1615);
   U2026 : INV3 port map( A => n1613, Q => n1010);
   U2027 : NAND22 port map( A => position1_n1323, B => n621, Q => n1614);
   U2028 : AOI211 port map( A => n1301, B => n515, C => n2013, Q => n2014);
   U2029 : AOI221 port map( A => n2012, B => n2011, C => n518, D => 
                           position1_n1547, Q => n2013);
   U2030 : AOI211 port map( A => n1082, B => n35, C => n1679, Q => n1680);
   U2031 : AOI221 port map( A => n1678, B => n1677, C => n518, D => 
                           position1_n1351, Q => n1679);
   U2032 : AOI221 port map( A => n2055, B => n2054, C => n625, D => n1307, Q =>
                           n2057);
   U2033 : INV3 port map( A => position1_N1556_port, Q => n1307);
   U2034 : NAND22 port map( A => position1_N1556_port, B => n246, Q => n2054);
   U2035 : AOI221 port map( A => position1_N1555_port, B => n67, C => n2053, D 
                           => n2052, Q => n2055);
   U2036 : AOI221 port map( A => n1721, B => n1720, C => n625, D => n1088, Q =>
                           n1723);
   U2037 : INV3 port map( A => position1_N1973, Q => n1088);
   U2038 : NAND22 port map( A => position1_N1973, B => n246, Q => n1720);
   U2039 : AOI221 port map( A => position1_N1972, B => n245, C => n1719, D => 
                           n1718, Q => n1721);
   U2040 : AOI221 port map( A => n1176, B => n282, C => n1874, D => n1873, Q =>
                           n1876);
   U2041 : NAND22 port map( A => n617, B => position1_n1469, Q => n1873);
   U2042 : AOI221 port map( A => n1872, B => n1871, C => n470, D => 
                           position1_n1470, Q => n1874);
   U2043 : NAND22 port map( A => n1177, B => n46, Q => n1871);
   U2044 : AOI221 port map( A => n957, B => n254, C => n1540, D => n1539, Q => 
                           n1542);
   U2045 : NAND22 port map( A => n617, B => position1_n1273, Q => n1539);
   U2046 : AOI221 port map( A => n1538, B => n1537, C => n471, D => 
                           position1_n1274, Q => n1540);
   U2047 : NAND22 port map( A => n958, B => n46, Q => n1537);
   U2048 : AOI221 port map( A => n2059, B => n2058, C => n622, D => n1309, Q =>
                           n2061);
   U2049 : INV3 port map( A => position1_N1558_port, Q => n1309);
   U2050 : NAND22 port map( A => position1_N1558_port, B => n250, Q => n2058);
   U2051 : AOI221 port map( A => position1_N1557_port, B => n248, C => n2057, D
                           => n2056, Q => n2059);
   U2052 : AOI221 port map( A => n1725, B => n1724, C => n622, D => n1090, Q =>
                           n1727);
   U2053 : INV3 port map( A => position1_N1975, Q => n1090);
   U2054 : NAND22 port map( A => position1_N1975, B => n250, Q => n1724);
   U2055 : AOI221 port map( A => position1_N1974, B => n42, C => n1723, D => 
                           n1722, Q => n1725);
   U2056 : AOI221 port map( A => n2063, B => n2062, C => n618, D => n1311, Q =>
                           n2065);
   U2057 : INV3 port map( A => position1_N1560_port, Q => n1311);
   U2058 : NAND22 port map( A => position1_N1560_port, B => n101, Q => n2062);
   U2059 : AOI221 port map( A => position1_N1559_port, B => n252, C => n2061, D
                           => n2060, Q => n2063);
   U2060 : AOI221 port map( A => n1729, B => n1728, C => n614, D => n1092, Q =>
                           n1731);
   U2061 : INV3 port map( A => position1_N1977, Q => n1092);
   U2062 : NAND22 port map( A => position1_N1977, B => n282, Q => n1728);
   U2063 : AOI221 port map( A => position1_N1976, B => n252, C => n1727, D => 
                           n1726, Q => n1729);
   U2064 : AOI221 port map( A => n2067, B => n2066, C => n613, D => n1313, Q =>
                           n2069);
   U2065 : INV3 port map( A => position1_N1562_port, Q => n1313);
   U2066 : NAND22 port map( A => position1_N1562_port, B => n286, Q => n2066);
   U2067 : AOI221 port map( A => position1_N1561_port, B => n256, C => n2065, D
                           => n2064, Q => n2067);
   U2068 : AOI221 port map( A => n1733, B => n1732, C => n612, D => n1094, Q =>
                           n1735);
   U2069 : INV3 port map( A => position1_N1979, Q => n1094);
   U2070 : NAND22 port map( A => position1_N1979, B => n286, Q => n1732);
   U2071 : AOI221 port map( A => position1_N1978, B => n284, C => n1731, D => 
                           n1730, Q => n1733);
   U2072 : AOI221 port map( A => n2071, B => n2070, C => n608, D => n1315, Q =>
                           n2073);
   U2073 : INV3 port map( A => position1_N1564_port, Q => n1315);
   U2074 : NAND22 port map( A => position1_N1564_port, B => n39, Q => n2070);
   U2075 : AOI221 port map( A => position1_N1563_port, B => n259, C => n2069, D
                           => n2068, Q => n2071);
   U2076 : AOI221 port map( A => n1737, B => n1736, C => n608, D => n1096, Q =>
                           n1739);
   U2077 : INV3 port map( A => position1_N1981, Q => n1096);
   U2078 : NAND22 port map( A => position1_N1981, B => n290, Q => n1736);
   U2079 : AOI221 port map( A => position1_N1980, B => n259, C => n1735, D => 
                           n1734, Q => n1737);
   U2080 : AOI221 port map( A => n2075, B => n2074, C => n604, D => n1317, Q =>
                           n2077);
   U2081 : INV3 port map( A => position1_N1566_port, Q => n1317);
   U2082 : NAND22 port map( A => position1_N1566_port, B => n40, Q => n2074);
   U2083 : AOI221 port map( A => position1_N1565_port, B => n263, C => n2073, D
                           => n2072, Q => n2075);
   U2084 : AOI221 port map( A => n1741, B => n1740, C => n604, D => n1098, Q =>
                           n1743);
   U2085 : INV3 port map( A => position1_N1983, Q => n1098);
   U2086 : NAND22 port map( A => position1_N1983, B => n294, Q => n1740);
   U2087 : AOI221 port map( A => position1_N1982, B => n44, C => n1739, D => 
                           n1738, Q => n1741);
   U2088 : AOI221 port map( A => n2079, B => n2078, C => n600, D => n1319, Q =>
                           n2081);
   U2089 : INV3 port map( A => position1_N1568_port, Q => n1319);
   U2090 : NAND22 port map( A => position1_N1568_port, B => n68, Q => n2078);
   U2091 : AOI221 port map( A => position1_N1567_port, B => n267, C => n2077, D
                           => n2076, Q => n2079);
   U2092 : AOI221 port map( A => n1745, B => n1744, C => n600, D => n1100, Q =>
                           n1747);
   U2093 : INV3 port map( A => position1_N1985, Q => n1100);
   U2094 : NAND22 port map( A => position1_N1985, B => n298, Q => n1744);
   U2095 : AOI221 port map( A => position1_N1984, B => n43, C => n1743, D => 
                           n1742, Q => n1745);
   U2096 : AOI221 port map( A => n1806, B => n1805, C => n608, D => 
                           position1_n1417, Q => n1808);
   U2097 : NAND22 port map( A => n1112, B => n261, Q => n1805);
   U2098 : AOI221 port map( A => n1114, B => n288, C => n1113, D => n1804, Q =>
                           n1806);
   U2099 : INV3 port map( A => position1_n1417, Q => n1112);
   U2100 : AOI221 port map( A => n1472, B => n1471, C => n608, D => 
                           position1_n1221, Q => n1474);
   U2101 : NAND22 port map( A => n893, B => n290, Q => n1471);
   U2102 : AOI221 port map( A => n895, B => n259, C => n894, D => n1470, Q => 
                           n1472);
   U2103 : INV3 port map( A => position1_n1221, Q => n893);
   U2104 : AOI221 port map( A => n1810, B => n1809, C => n604, D => 
                           position1_n1415, Q => n1812);
   U2105 : NAND22 port map( A => n1110, B => n294, Q => n1809);
   U2106 : AOI221 port map( A => n1111, B => n44, C => n1808, D => n1807, Q => 
                           n1810);
   U2107 : INV3 port map( A => position1_n1415, Q => n1110);
   U2108 : AOI221 port map( A => n1476, B => n1475, C => n604, D => 
                           position1_n1219, Q => n1478);
   U2109 : NAND22 port map( A => n891, B => n265, Q => n1475);
   U2110 : AOI221 port map( A => n892, B => n263, C => n1474, D => n1473, Q => 
                           n1476);
   U2111 : INV3 port map( A => position1_n1219, Q => n891);
   U2112 : AOI221 port map( A => n1814, B => n1813, C => n600, D => 
                           position1_n1413, Q => n1816);
   U2113 : NAND22 port map( A => n1108, B => n269, Q => n1813);
   U2114 : AOI221 port map( A => n1109, B => n43, C => n1812, D => n1811, Q => 
                           n1814);
   U2115 : INV3 port map( A => position1_n1413, Q => n1108);
   U2116 : AOI221 port map( A => n1480, B => n1479, C => n600, D => 
                           position1_n1217, Q => n1482);
   U2117 : NAND22 port map( A => n889, B => n298, Q => n1479);
   U2118 : AOI221 port map( A => n890, B => n267, C => n1478, D => n1477, Q => 
                           n1480);
   U2119 : INV3 port map( A => position1_n1217, Q => n889);
   U2120 : AOI221 port map( A => n1180, B => n274, C => n1866, D => n1865, Q =>
                           n1868);
   U2121 : NAND22 port map( A => n624, B => position1_n1473, Q => n1865);
   U2122 : AOI221 port map( A => n1864, B => n1863, C => n629, D => 
                           position1_n1474, Q => n1866);
   U2123 : NAND22 port map( A => n1181, B => n67, Q => n1863);
   U2124 : AOI221 port map( A => n961, B => n274, C => n1532, D => n1531, Q => 
                           n1534);
   U2125 : NAND22 port map( A => n625, B => position1_n1277, Q => n1531);
   U2126 : AOI221 port map( A => n1530, B => n1529, C => n629, D => 
                           position1_n1278, Q => n1532);
   U2127 : NAND22 port map( A => n962, B => n272, Q => n1529);
   U2128 : AOI221 port map( A => n1178, B => n278, C => n1870, D => n1869, Q =>
                           n1872);
   U2129 : NAND22 port map( A => n622, B => position1_n1471, Q => n1869);
   U2130 : AOI221 port map( A => n1868, B => n1867, C => n469, D => 
                           position1_n1472, Q => n1870);
   U2131 : NAND22 port map( A => n1179, B => n42, Q => n1867);
   U2132 : AOI221 port map( A => n959, B => n250, C => n1536, D => n1535, Q => 
                           n1538);
   U2133 : NAND22 port map( A => n622, B => position1_n1275, Q => n1535);
   U2134 : AOI221 port map( A => n1534, B => n1533, C => position1_N2457, D => 
                           position1_n1276, Q => n1536);
   U2135 : NAND22 port map( A => n960, B => n248, Q => n1533);
   U2136 : AOI221 port map( A => n1172, B => n261, C => n1882, D => n1881, Q =>
                           n1884);
   U2137 : NAND22 port map( A => n607, B => position1_n1465, Q => n1881);
   U2138 : AOI221 port map( A => n1880, B => n1879, C => n474, D => 
                           position1_n1466, Q => n1882);
   U2139 : NAND22 port map( A => n1173, B => n47, Q => n1879);
   U2140 : AOI221 port map( A => n953, B => n290, C => n1548, D => n1547, Q => 
                           n1550);
   U2141 : NAND22 port map( A => n607, B => position1_n1269, Q => n1547);
   U2142 : AOI221 port map( A => n1546, B => n1545, C => n474, D => 
                           position1_n1270, Q => n1548);
   U2143 : NAND22 port map( A => n954, B => n47, Q => n1545);
   U2144 : AOI221 port map( A => n1170, B => n294, C => n1886, D => n1885, Q =>
                           n1888);
   U2145 : NAND22 port map( A => n603, B => position1_n1463, Q => n1885);
   U2146 : AOI221 port map( A => n1884, B => n1883, C => n475, D => 
                           position1_n1464, Q => n1886);
   U2147 : NAND22 port map( A => n1171, B => n44, Q => n1883);
   U2148 : AOI221 port map( A => n951, B => n265, C => n1552, D => n1551, Q => 
                           n1554);
   U2149 : NAND22 port map( A => n603, B => position1_n1267, Q => n1551);
   U2150 : AOI221 port map( A => n1550, B => n1549, C => position1_N2449, D => 
                           position1_n1268, Q => n1552);
   U2151 : NAND22 port map( A => n952, B => n44, Q => n1549);
   U2152 : AOI221 port map( A => n1182, B => n273, C => n1862, D => n1861, Q =>
                           n1864);
   U2153 : NAND22 port map( A => n633, B => position1_n1475, Q => n1861);
   U2154 : AOI211 port map( A => n519, B => position1_n1476, C => n1860, Q => 
                           n1862);
   U2155 : AOI2111 port map( A => n1183, B => n35, C => n1184, D => n1185, Q =>
                           n1860);
   U2156 : AOI221 port map( A => n963, B => n273, C => n1528, D => n1527, Q => 
                           n1530);
   U2157 : NAND22 port map( A => n633, B => position1_n1279, Q => n1527);
   U2158 : AOI211 port map( A => n519, B => position1_n1280, C => n1526, Q => 
                           n1528);
   U2159 : AOI2111 port map( A => n964, B => n35, C => n965, D => n966, Q => 
                           n1526);
   U2160 : AOI221 port map( A => n1174, B => n286, C => n1878, D => n1877, Q =>
                           n1880);
   U2161 : NAND22 port map( A => n612, B => position1_n1467, Q => n1877);
   U2162 : AOI221 port map( A => n1876, B => n1875, C => n472, D => 
                           position1_n1468, Q => n1878);
   U2163 : NAND22 port map( A => n1175, B => n41, Q => n1875);
   U2164 : AOI221 port map( A => n955, B => n286, C => n1544, D => n1543, Q => 
                           n1546);
   U2165 : NAND22 port map( A => n612, B => position1_n1271, Q => n1543);
   U2166 : AOI221 port map( A => n1542, B => n1541, C => position1_N2453, D => 
                           position1_n1272, Q => n1544);
   U2167 : NAND22 port map( A => n956, B => n256, Q => n1541);
   U2168 : AOI221 port map( A => n1790, B => n1789, C => n625, D => 
                           position1_n1425, Q => n1792);
   U2169 : NAND22 port map( A => n1121, B => n274, Q => n1789);
   U2170 : AOI221 port map( A => n1122, B => n272, C => n1788, D => n1787, Q =>
                           n1790);
   U2171 : INV3 port map( A => position1_n1425, Q => n1121);
   U2172 : AOI221 port map( A => n1456, B => n1455, C => n625, D => 
                           position1_n1229, Q => n1458);
   U2173 : NAND22 port map( A => n902, B => n246, Q => n1455);
   U2174 : AOI221 port map( A => n903, B => n245, C => n1454, D => n1453, Q => 
                           n1456);
   U2175 : INV3 port map( A => position1_n1229, Q => n902);
   U2176 : AOI221 port map( A => n1794, B => n1793, C => n622, D => 
                           position1_n1423, Q => n1796);
   U2177 : NAND22 port map( A => n1119, B => n278, Q => n1793);
   U2178 : AOI221 port map( A => n1120, B => n276, C => n1792, D => n1791, Q =>
                           n1794);
   U2179 : INV3 port map( A => position1_n1423, Q => n1119);
   U2180 : AOI221 port map( A => n1460, B => n1459, C => n622, D => 
                           position1_n1227, Q => n1462);
   U2181 : NAND22 port map( A => n900, B => n250, Q => n1459);
   U2182 : AOI221 port map( A => n901, B => n248, C => n1458, D => n1457, Q => 
                           n1460);
   U2183 : INV3 port map( A => position1_n1227, Q => n900);
   U2184 : AOI221 port map( A => n2051, B => n2050, C => n634, D => n1305, Q =>
                           n2053);
   U2185 : INV3 port map( A => position1_N1554_port, Q => n1305);
   U2186 : NAND22 port map( A => position1_N1554_port, B => n630, Q => n2050);
   U2187 : AOI211 port map( A => position1_N1553_port, B => n515, C => n2049, Q
                           => n2051);
   U2188 : AOI221 port map( A => n1717, B => n1716, C => n634, D => n1086, Q =>
                           n1719);
   U2189 : INV3 port map( A => position1_N1971, Q => n1086);
   U2190 : NAND22 port map( A => position1_N1971, B => n273, Q => n1716);
   U2191 : AOI211 port map( A => position1_N1970, B => n35, C => n1715, Q => 
                           n1717);
   U2192 : INV3 port map( A => position1_N1656, Q => n1265);
   U2193 : AOI211 port map( A => position1_N1655, B => n515, C => n1974, Q => 
                           n1975);
   U2194 : AOI221 port map( A => n1973, B => n1972, C => n518, D => n1266, Q =>
                           n1974);
   U2195 : INV3 port map( A => position1_N2073, Q => n1046);
   U2196 : AOI211 port map( A => position1_N2072, B => n35, C => n1640, Q => 
                           n1641);
   U2197 : AOI221 port map( A => n1639, B => n1638, C => n518, D => n1047, Q =>
                           n1640);
   U2198 : INV3 port map( A => n167, Q => position1_sub_216_I2_carry_8_port);
   U2199 : NOR21 port map( A => n515, B => position1_N1553_port, Q => n167);
   U2200 : INV3 port map( A => n173, Q => position1_sub_226_I2_carry_8_port);
   U2201 : NOR21 port map( A => n515, B => position1_N1970, Q => n173);
   U2202 : INV3 port map( A => position1_N1519_port, Q => n523);
   U2203 : INV3 port map( A => position1_N1936, Q => n557);
   U2204 : AOI211 port map( A => n634, B => n1786, C => n1123, Q => n1788);
   U2205 : INV3 port map( A => n1785, Q => n1123);
   U2206 : NAND22 port map( A => n1124, B => n35, Q => n1786);
   U2207 : AOI211 port map( A => n634, B => n1452, C => n904, Q => n1454);
   U2208 : INV3 port map( A => n1451, Q => n904);
   U2209 : NAND22 port map( A => n905, B => n35, Q => n1452);
   U2210 : NAND22 port map( A => position1_n1545, B => n627, Q => n2010);
   U2211 : NAND22 port map( A => position1_n1349, B => n627, Q => n1676);
   U2212 : NAND22 port map( A => position1_n1544, B => n624, Q => n2020);
   U2213 : NAND22 port map( A => position1_n1348, B => n624, Q => n1686);
   U2214 : NOR21 port map( A => n620, B => position1_n1519, Q => n1946);
   U2215 : NOR21 port map( A => n621, B => position1_n1323, Q => n1612);
   U2216 : BUF2 port map( A => position1_n1152, Q => n487);
   U2217 : NAND22 port map( A => n596, B => position1_n1460, Q => n1894);
   U2218 : NAND22 port map( A => n595, B => position1_n1264, Q => n1560);
   U2219 : NOR21 port map( A => n52, B => n632, Q => n2086);
   U2220 : NOR21 port map( A => n51, B => n632, Q => n1752);
   U2221 : BUF2 port map( A => n102, Q => n591);
   U2222 : BUF2 port map( A => n592, Q => n590);
   U2223 : NAND22 port map( A => n612, B => position1_n1419, Q => n1804);
   U2224 : NAND22 port map( A => n612, B => position1_n1223, Q => n1470);
   U2225 : NAND22 port map( A => position1_N2449, B => position1_n1416, Q => 
                           n1807);
   U2226 : NAND22 port map( A => position1_N2449, B => position1_n1220, Q => 
                           n1473);
   U2227 : NAND22 port map( A => position1_N2447, B => position1_n1414, Q => 
                           n1811);
   U2228 : NAND22 port map( A => position1_N2447, B => position1_n1218, Q => 
                           n1477);
   U2229 : NAND22 port map( A => n595, B => position1_n1412, Q => n1815);
   U2230 : NAND22 port map( A => n596, B => position1_n1216, Q => n1481);
   U2231 : NAND22 port map( A => n629, B => position1_n1426, Q => n1787);
   U2232 : NAND22 port map( A => n629, B => position1_n1230, Q => n1453);
   U2233 : NAND22 port map( A => position1_N2457, B => position1_n1424, Q => 
                           n1791);
   U2234 : NAND22 port map( A => position1_N2457, B => position1_n1228, Q => 
                           n1457);
   U2235 : NAND22 port map( A => n471, B => position1_n1422, Q => n1795);
   U2236 : NAND22 port map( A => n471, B => position1_n1226, Q => n1461);
   U2237 : NAND22 port map( A => position1_n1445, B => n616, Q => n1839);
   U2238 : NAND22 port map( A => position1_n1249, B => n616, Q => n1505);
   U2239 : NAND22 port map( A => position1_n1531, B => n594, Q => n2044);
   U2240 : NAND22 port map( A => position1_n1335, B => n594, Q => n1710);
   U2241 : NOR21 port map( A => n602, B => position1_n1487, Q => n1926);
   U2242 : NOR21 port map( A => n602, B => position1_n1291, Q => n1592);
   U2243 : NOR21 port map( A => n624, B => n1263, Q => n1980);
   U2244 : INV3 port map( A => position1_N1658, Q => n1263);
   U2245 : NOR21 port map( A => n623, B => n1044, Q => n1646);
   U2246 : INV3 port map( A => position1_N2075, Q => n1044);
   U2247 : NOR21 port map( A => n615, B => n1259, Q => n1988);
   U2248 : INV3 port map( A => position1_N1662, Q => n1259);
   U2249 : NOR21 port map( A => n616, B => n1040, Q => n1654);
   U2250 : INV3 port map( A => position1_N2079, Q => n1040);
   U2251 : NOR21 port map( A => n610, B => n1257, Q => n1992);
   U2252 : INV3 port map( A => position1_N1664, Q => n1257);
   U2253 : NOR21 port map( A => n610, B => n1038, Q => n1658);
   U2254 : INV3 port map( A => position1_N2081, Q => n1038);
   U2255 : NOR21 port map( A => n606, B => n1255, Q => n1996);
   U2256 : INV3 port map( A => position1_N1666, Q => n1255);
   U2257 : NOR21 port map( A => n606, B => n1036, Q => n1662);
   U2258 : INV3 port map( A => position1_N2083, Q => n1036);
   U2259 : NOR21 port map( A => n602, B => n1253, Q => n2000);
   U2260 : INV3 port map( A => position1_N1668, Q => n1253);
   U2261 : NOR21 port map( A => n602, B => n1034, Q => n1666);
   U2262 : INV3 port map( A => position1_N2085, Q => n1034);
   U2263 : NOR21 port map( A => n598, B => n1251, Q => n2004);
   U2264 : INV3 port map( A => position1_N1670, Q => n1251);
   U2265 : NOR21 port map( A => n598, B => n1032, Q => n1670);
   U2266 : INV3 port map( A => position1_N2087, Q => n1032);
   U2267 : NOR21 port map( A => n620, B => n1261, Q => n1984);
   U2268 : INV3 port map( A => position1_N1660, Q => n1261);
   U2269 : NOR21 port map( A => n620, B => n1042, Q => n1650);
   U2270 : INV3 port map( A => position1_N2077, Q => n1042);
   U2271 : NAND22 port map( A => n629, B => n1306, Q => n2052);
   U2272 : INV3 port map( A => position1_N1555_port, Q => n1306);
   U2273 : NAND22 port map( A => n628, B => n1087, Q => n1718);
   U2274 : INV3 port map( A => position1_N1972, Q => n1087);
   U2275 : NAND22 port map( A => n469, B => n1308, Q => n2056);
   U2276 : INV3 port map( A => position1_N1557_port, Q => n1308);
   U2277 : NAND22 port map( A => n469, B => n1089, Q => n1722);
   U2278 : INV3 port map( A => position1_N1974, Q => n1089);
   U2279 : NAND22 port map( A => n470, B => n1310, Q => n2060);
   U2280 : INV3 port map( A => position1_N1559_port, Q => n1310);
   U2281 : NAND22 port map( A => n470, B => n1091, Q => n1726);
   U2282 : INV3 port map( A => position1_N1976, Q => n1091);
   U2283 : NAND22 port map( A => n472, B => n1312, Q => n2064);
   U2284 : INV3 port map( A => position1_N1561_port, Q => n1312);
   U2285 : NAND22 port map( A => n472, B => n1093, Q => n1730);
   U2286 : INV3 port map( A => position1_N1978, Q => n1093);
   U2287 : NAND22 port map( A => n474, B => n1314, Q => n2068);
   U2288 : INV3 port map( A => position1_N1563_port, Q => n1314);
   U2289 : NAND22 port map( A => n474, B => n1095, Q => n1734);
   U2290 : INV3 port map( A => position1_N1980, Q => n1095);
   U2291 : NAND22 port map( A => n475, B => n1316, Q => n2072);
   U2292 : INV3 port map( A => position1_N1565_port, Q => n1316);
   U2293 : NAND22 port map( A => n475, B => n1097, Q => n1738);
   U2294 : INV3 port map( A => position1_N1982, Q => n1097);
   U2295 : NAND22 port map( A => n476, B => n1318, Q => n2076);
   U2296 : INV3 port map( A => position1_N1567_port, Q => n1318);
   U2297 : NAND22 port map( A => n476, B => n1099, Q => n1742);
   U2298 : INV3 port map( A => position1_N1984, Q => n1099);
   U2299 : INV3 port map( A => n1846, Q => n1143);
   U2300 : AOI2111 port map( A => n1144, B => n47, C => n1845, D => n1844, Q =>
                           n1846);
   U2301 : NOR21 port map( A => n610, B => position1_n1443, Q => n1845);
   U2302 : AOI2111 port map( A => n611, B => position1_n1443, C => n1843, D => 
                           n1842, Q => n1844);
   U2303 : INV3 port map( A => n1512, Q => n924);
   U2304 : AOI2111 port map( A => n925, B => n259, C => n1511, D => n1510, Q =>
                           n1512);
   U2305 : NOR21 port map( A => n610, B => position1_n1247, Q => n1511);
   U2306 : AOI2111 port map( A => n611, B => position1_n1247, C => n1509, D => 
                           n1508, Q => n1510);
   U2307 : INV3 port map( A => n1929, Q => n1195);
   U2308 : NOR21 port map( A => n1196, B => n43, Q => n1928);
   U2309 : INV3 port map( A => n1595, Q => n976);
   U2310 : NOR21 port map( A => n977, B => n267, Q => n1594);
   U2311 : INV3 port map( A => n1799, Q => n1116);
   U2312 : AOI221 port map( A => n1798, B => n1797, C => n618, D => 
                           position1_n1421, Q => n1799);
   U2313 : NAND22 port map( A => n1117, B => n254, Q => n1797);
   U2314 : AOI221 port map( A => n1118, B => n46, C => n1796, D => n1795, Q => 
                           n1798);
   U2315 : INV3 port map( A => n1465, Q => n897);
   U2316 : AOI221 port map( A => n1464, B => n1463, C => n618, D => 
                           position1_n1225, Q => n1465);
   U2317 : NAND22 port map( A => n898, B => n282, Q => n1463);
   U2318 : AOI221 port map( A => n899, B => n252, C => n1462, D => n1461, Q => 
                           n1464);
   U2319 : INV3 port map( A => n1803, Q => n1113);
   U2320 : NOR21 port map( A => position1_n1419, B => n611, Q => n1801);
   U2321 : INV3 port map( A => n1469, Q => n894);
   U2322 : NOR21 port map( A => position1_n1223, B => n611, Q => n1467);
   U2323 : INV3 port map( A => n2090, Q => n1344);
   U2324 : NOR21 port map( A => n66, B => n624, Q => n2090);
   U2325 : INV3 port map( A => n1756, Q => n1343);
   U2326 : NOR21 port map( A => n59, B => n624, Q => n1756);
   U2327 : INV3 port map( A => n2094, Q => n1340);
   U2328 : NOR21 port map( A => n65, B => n621, Q => n2094);
   U2329 : INV3 port map( A => n1760, Q => n1339);
   U2330 : NOR21 port map( A => n58, B => n621, Q => n1760);
   U2331 : INV3 port map( A => n2098, Q => n1336);
   U2332 : NOR21 port map( A => n64, B => n616, Q => n2098);
   U2333 : INV3 port map( A => n1764, Q => n1335);
   U2334 : NOR21 port map( A => n57, B => n617, Q => n1764);
   U2335 : INV3 port map( A => n2102, Q => n1332);
   U2336 : NOR21 port map( A => n63, B => n611, Q => n2102);
   U2337 : INV3 port map( A => n1768, Q => n1331);
   U2338 : NOR21 port map( A => n56, B => n611, Q => n1768);
   U2339 : INV3 port map( A => n2106, Q => n1328);
   U2340 : NOR21 port map( A => n62, B => n607, Q => n2106);
   U2341 : INV3 port map( A => n1772, Q => n1327);
   U2342 : NOR21 port map( A => n55, B => n607, Q => n1772);
   U2343 : INV3 port map( A => n2110, Q => n1324);
   U2344 : NOR21 port map( A => n61, B => n603, Q => n2110);
   U2345 : INV3 port map( A => n1776, Q => n1323);
   U2346 : NOR21 port map( A => n54, B => n603, Q => n1776);
   U2347 : INV3 port map( A => n2114, Q => n1320);
   U2348 : NOR21 port map( A => n60, B => n599, Q => n2114);
   U2349 : INV3 port map( A => n1780, Q => n1101);
   U2350 : NOR21 port map( A => n53, B => n599, Q => n1780);
   U2351 : INV3 port map( A => n1898, Q => n1186);
   U2352 : NOR21 port map( A => n598, B => position1_n1485, Q => n1898);
   U2353 : INV3 port map( A => n1564, Q => n967);
   U2354 : NOR21 port map( A => n598, B => position1_n1289, Q => n1564);
   U2355 : INV3 port map( A => n1800, Q => n1115);
   U2356 : NAND22 port map( A => position1_N2453, B => position1_n1420, Q => 
                           n1800);
   U2357 : INV3 port map( A => n1466, Q => n896);
   U2358 : NAND22 port map( A => position1_N2453, B => position1_n1224, Q => 
                           n1466);
   U2359 : BUF2 port map( A => n102, Q => n592);
   U2360 : NOR40 port map( A => n818, B => n827, C => gensync1_N167, D => 
                           gensync1_N168, Q => gensync1_N129);
   U2361 : INV3 port map( A => n1373, Q => n827);
   U2362 : INV3 port map( A => n1372, Q => n818);
   U2363 : NOR31 port map( A => gensync1_N166, B => gensync1_comptY_9_port, C 
                           => gensync1_N165, Q => n1373);
   U2364 : NOR40 port map( A => gensync1_N169, B => gensync1_N170, C => 
                           gensync1_N171, D => gensync1_N172, Q => n1372);
   U2365 : AOI2111 port map( A => gensync1_N176, B => n872, C => gensync1_N174,
                           D => n477, Q => gensync1_N69);
   U2366 : INV3 port map( A => n1383, Q => n872);
   U2367 : NOR40 port map( A => gensync1_N177, B => gensync1_N178, C => 
                           gensync1_N179, D => n873, Q => n1383);
   U2368 : INV3 port map( A => n1382, Q => n873);
   U2369 : AOI211 port map( A => n477, B => n1381, C => gensync1_N174, Q => 
                           gensync1_N72);
   U2370 : NAND31 port map( A => n1380, B => n7, C => n1379, Q => n1381);
   U2371 : NOR31 port map( A => gensync1_N178, B => gensync1_N176, C => 
                           gensync1_N177, Q => n1379);
   U2372 : NAND22 port map( A => n816, B => n3, Q => gensync1_n99);
   U2373 : NAND41 port map( A => position1_n860, B => position1_n861, C => 
                           position1_n862, D => position1_n863, Q => 
                           position1_n1587);
   U2374 : NAND22 port map( A => position1_y_sum_23_port, B => n512, Q => 
                           position1_n861);
   U2375 : NAND22 port map( A => position1_N1225_port, B => n640, Q => 
                           position1_n863);
   U2376 : AOI221 port map( A => position1_N558, B => n514, C => 
                           position1_N1002_port, D => n643, Q => position1_n862
                           );
   U2377 : NAND41 port map( A => position1_n960, B => position1_n961, C => 
                           position1_n962, D => position1_n963, Q => 
                           position1_n1612);
   U2378 : NAND22 port map( A => position1_x_sum_23_port, B => n510, Q => 
                           position1_n961);
   U2379 : NAND22 port map( A => position1_N1200_port, B => n637, Q => 
                           position1_n963);
   U2380 : AOI221 port map( A => position1_N508, B => n513, C => 
                           position1_N927_port, D => n641, Q => position1_n962)
                           ;
   U2381 : NAND41 port map( A => position1_n964, B => position1_n965, C => 
                           position1_n966, D => position1_n967, Q => 
                           position1_n1613);
   U2382 : NAND22 port map( A => position1_x_sum_22_port, B => n510, Q => 
                           position1_n965);
   U2383 : NAND22 port map( A => position1_N1199_port, B => n637, Q => 
                           position1_n967);
   U2384 : AOI221 port map( A => position1_N507, B => n513, C => 
                           position1_N926_port, D => n641, Q => position1_n966)
                           ;
   U2385 : NAND41 port map( A => position1_n852, B => position1_n853, C => 
                           position1_n854, D => position1_n855, Q => 
                           position1_n1586);
   U2386 : NAND22 port map( A => position1_y_sum_24_port, B => n512, Q => 
                           position1_n853);
   U2387 : NAND22 port map( A => position1_N1226_port, B => n640, Q => 
                           position1_n855);
   U2388 : AOI221 port map( A => position1_N559, B => n514, C => 
                           position1_N1003_port, D => n643, Q => position1_n854
                           );
   U2389 : NAND41 port map( A => position1_n956, B => position1_n957, C => 
                           position1_n958, D => position1_n959, Q => 
                           position1_n1611);
   U2390 : NAND22 port map( A => position1_x_sum_24_port, B => n675, Q => 
                           position1_n957);
   U2391 : NAND22 port map( A => position1_N1201_port, B => n638, Q => 
                           position1_n959);
   U2392 : AOI221 port map( A => position1_N509, B => n513, C => 
                           position1_N928_port, D => n641, Q => position1_n958)
                           ;
   U2393 : NOR31 port map( A => n1366, B => n1365, C => n1364, Q => n1367);
   U2394 : NAND22 port map( A => gensync1_N170, B => gensync1_N168, Q => n1364)
                           ;
   U2395 : NAND31 port map( A => gensync1_N165, B => gensync1_N166, C => 
                           gensync1_N169, Q => n1365);
   U2396 : NAND41 port map( A => gensync1_N173, B => gensync1_N171, C => 
                           gensync1_N172, D => gensync1_N167, Q => n1366);
   U2397 : NOR40 port map( A => n1371, B => gensync1_N166, C => 
                           gensync1_comptY_9_port, D => gensync1_N165, Q => 
                           gensync1_N132);
   U2398 : NOR21 port map( A => gensync1_N167, B => gensync1_N168, Q => n1368);
   U2399 : NAND22 port map( A => gensync1_N169, B => gensync1_N170, Q => n1369)
                           ;
   U2400 : INV3 port map( A => gensync1_n98, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port);
   U2401 : NAND22 port map( A => n816, B => gensync1_N138, Q => gensync1_n98);
   U2402 : XOR21 port map( A => gensync1_N173, B => gensync1_N172, Q => 
                           gensync1_N138);
   U2403 : NAND31 port map( A => gensync1_N172, B => gensync1_N173, C => 
                           gensync1_N171, Q => n1370);
   U2404 : NOR21 port map( A => n199, B => n76, Q => 
                           position1_r409_carry_13_port);
   U2405 : INV3 port map( A => position1_r409_carry_12_port, Q => n199);
   U2406 : NOR21 port map( A => n183, B => n82, Q => 
                           position1_r406_carry_13_port);
   U2407 : INV3 port map( A => position1_r406_carry_12_port, Q => n183);
   U2408 : NOR21 port map( A => n197, B => n69, Q => 
                           position1_r409_carry_11_port);
   U2409 : INV3 port map( A => position1_r409_carry_10_port, Q => n197);
   U2410 : NOR21 port map( A => n181, B => n70, Q => 
                           position1_r406_carry_11_port);
   U2411 : INV3 port map( A => position1_r406_carry_10_port, Q => n181);
   U2412 : NOR21 port map( A => n196, B => n51, Q => 
                           position1_r409_carry_10_port);
   U2413 : INV3 port map( A => position1_r409_carry_9_port, Q => n196);
   U2414 : NOR21 port map( A => n180, B => n52, Q => 
                           position1_r406_carry_10_port);
   U2415 : INV3 port map( A => position1_r406_carry_9_port, Q => n180);
   U2416 : NOR21 port map( A => n198, B => n59, Q => 
                           position1_r409_carry_12_port);
   U2417 : INV3 port map( A => position1_r409_carry_11_port, Q => n198);
   U2418 : NOR21 port map( A => n182, B => n66, Q => 
                           position1_r406_carry_12_port);
   U2419 : INV3 port map( A => position1_r406_carry_11_port, Q => n182);
   U2420 : INV3 port map( A => gensync1_N66, Q => n874);
   U2421 : NOR40 port map( A => gensync1_N174, B => n477, C => gensync1_N176, D
                           => n1385, Q => gensync1_N66);
   U2422 : NOR21 port map( A => n1384, B => n6, Q => n1385);
   U2423 : AOI311 port map( A => gensync1_N180, B => gensync1_N181, C => 
                           gensync1_N179, D => gensync1_N178, Q => n1384);
   U2424 : NOR21 port map( A => n179, B => n98, Q => 
                           position1_r406_carry_1_port);
   U2425 : INV3 port map( A => n505, Q => n179);
   U2426 : AOI221 port map( A => position1_N428, B => n646, C => position1_N655
                           , D => n649, Q => position1_n860);
   U2427 : XOR21 port map( A => position1_y_sum_23_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_23_port, Q 
                           => position1_N655);
   U2428 : XOR21 port map( A => position1_N378, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_23_port, Q 
                           => position1_N428);
   U2429 : AOI221 port map( A => position1_N353_port, B => n644, C => 
                           position1_N630, D => n648, Q => position1_n960);
   U2430 : XOR21 port map( A => position1_x_sum_23_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_23_port, Q 
                           => position1_N630);
   U2431 : XOR21 port map( A => position1_N303, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_23_port, Q 
                           => position1_N353_port);
   U2432 : AOI221 port map( A => position1_N352_port, B => n644, C => 
                           position1_N629, D => n648, Q => position1_n964);
   U2433 : XOR21 port map( A => position1_x_sum_22_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_22_port, Q 
                           => position1_N629);
   U2434 : XOR21 port map( A => position1_N302, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_22_port, Q 
                           => position1_N352_port);
   U2435 : AOI221 port map( A => position1_N429, B => n646, C => position1_N656
                           , D => n649, Q => position1_n852);
   U2436 : XOR21 port map( A => 
                           position1_dp_cluster_5_add_179_aco_carry_24_port, B 
                           => position1_y_sum_24_port, Q => position1_N656);
   U2437 : XOR21 port map( A => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_24_port, B 
                           => position1_N379, Q => position1_N429);
   U2438 : NOR21 port map( A => n410, B => n53, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_24_port);
   U2439 : AOI221 port map( A => position1_N354, B => n644, C => position1_N631
                           , D => n648, Q => position1_n956);
   U2440 : XOR21 port map( A => 
                           position1_dp_cluster_4_add_178_aco_carry_24_port, B 
                           => position1_x_sum_24_port, Q => position1_N631);
   U2441 : XOR21 port map( A => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_24_port, B 
                           => position1_N304, Q => position1_N354);
   U2442 : NOR21 port map( A => n395, B => n60, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_24_port);
   U2443 : INV3 port map( A => gensync1_n105, Q => n816);
   U2444 : NAND22 port map( A => gensync1_n106, B => gensync1_N135, Q => 
                           gensync1_n105);
   U2445 : NOR21 port map( A => gensync1_comptY_9_port, B => n1367, Q => 
                           gensync1_N135);
   U2446 : NOR21 port map( A => gensync1_N132, B => gensync1_N129, Q => 
                           gensync1_n106);
   U2447 : NOR21 port map( A => n507, B => n10, Q => n2135);
   U2448 : NOR21 port map( A => n507, B => n1, Q => n2136);
   U2449 : NOR21 port map( A => n195, B => n97, Q => 
                           position1_r409_carry_1_port);
   U2450 : INV3 port map( A => cam_y_0_port, Q => n195);
   U2451 : NOR21 port map( A => n200, B => n58, Q => 
                           position1_r409_carry_14_port);
   U2452 : INV3 port map( A => position1_r409_carry_13_port, Q => n200);
   U2453 : NOR21 port map( A => n184, B => n65, Q => 
                           position1_r406_carry_14_port);
   U2454 : INV3 port map( A => position1_r406_carry_13_port, Q => n184);
   U2455 : NOR21 port map( A => n202, B => n57, Q => 
                           position1_r409_carry_16_port);
   U2456 : INV3 port map( A => position1_r409_carry_15_port, Q => n202);
   U2457 : NOR21 port map( A => n186, B => n64, Q => 
                           position1_r406_carry_16_port);
   U2458 : INV3 port map( A => position1_r406_carry_15_port, Q => n186);
   U2459 : NOR21 port map( A => n204, B => n56, Q => 
                           position1_r409_carry_18_port);
   U2460 : INV3 port map( A => position1_r409_carry_17_port, Q => n204);
   U2461 : NOR21 port map( A => n188, B => n63, Q => 
                           position1_r406_carry_18_port);
   U2462 : INV3 port map( A => position1_r406_carry_17_port, Q => n188);
   U2463 : NOR21 port map( A => n206, B => n55, Q => 
                           position1_r409_carry_20_port);
   U2464 : INV3 port map( A => position1_r409_carry_19_port, Q => n206);
   U2465 : NOR21 port map( A => n190, B => n62, Q => 
                           position1_r406_carry_20_port);
   U2466 : INV3 port map( A => position1_r406_carry_19_port, Q => n190);
   U2467 : NOR21 port map( A => n208, B => n54, Q => 
                           position1_r409_carry_22_port);
   U2468 : INV3 port map( A => position1_r409_carry_21_port, Q => n208);
   U2469 : NOR21 port map( A => n192, B => n61, Q => 
                           position1_r406_carry_22_port);
   U2470 : INV3 port map( A => position1_r406_carry_21_port, Q => n192);
   U2471 : XOR21 port map( A => position1_r406_carry_24_port, B => 
                           position1_x_sum_24_port, Q => position1_N304);
   U2472 : NOR21 port map( A => n194, B => n60, Q => 
                           position1_r406_carry_24_port);
   U2473 : INV3 port map( A => position1_r406_carry_23_port, Q => n194);
   U2474 : NOR21 port map( A => n201, B => n75, Q => 
                           position1_r409_carry_15_port);
   U2475 : INV3 port map( A => position1_r409_carry_14_port, Q => n201);
   U2476 : NOR21 port map( A => n185, B => n81, Q => 
                           position1_r406_carry_15_port);
   U2477 : INV3 port map( A => position1_r406_carry_14_port, Q => n185);
   U2478 : NOR21 port map( A => n203, B => n74, Q => 
                           position1_r409_carry_17_port);
   U2479 : INV3 port map( A => position1_r409_carry_16_port, Q => n203);
   U2480 : NOR21 port map( A => n187, B => n80, Q => 
                           position1_r406_carry_17_port);
   U2481 : INV3 port map( A => position1_r406_carry_16_port, Q => n187);
   U2482 : NOR21 port map( A => n205, B => n73, Q => 
                           position1_r409_carry_19_port);
   U2483 : INV3 port map( A => position1_r409_carry_18_port, Q => n205);
   U2484 : NOR21 port map( A => n189, B => n79, Q => 
                           position1_r406_carry_19_port);
   U2485 : INV3 port map( A => position1_r406_carry_18_port, Q => n189);
   U2486 : NOR21 port map( A => n207, B => n72, Q => 
                           position1_r409_carry_21_port);
   U2487 : INV3 port map( A => position1_r409_carry_20_port, Q => n207);
   U2488 : NOR21 port map( A => n191, B => n78, Q => 
                           position1_r406_carry_21_port);
   U2489 : INV3 port map( A => position1_r406_carry_20_port, Q => n191);
   U2490 : NOR21 port map( A => n209, B => n71, Q => 
                           position1_r409_carry_23_port);
   U2491 : INV3 port map( A => position1_r409_carry_22_port, Q => n209);
   U2492 : NOR21 port map( A => n193, B => n77, Q => 
                           position1_r406_carry_23_port);
   U2493 : INV3 port map( A => position1_r406_carry_22_port, Q => n193);
   U2494 : XOR21 port map( A => position1_N1938, B => cam_y_0_port, Q => 
                           position1_N355);
   U2495 : XOR21 port map( A => position1_N1521_port, B => n505, Q => 
                           position1_N280);
   U2496 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_8_port, Q 
                           => n779);
   U2497 : NAND22 port map( A => n1363, B => position1_dp_cluster_6_N389, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_8_port);
   U2498 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_8_port, Q 
                           => n869);
   U2499 : NAND22 port map( A => n1363, B => position1_dp_cluster_7_N314, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_8_port);
   U2500 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_8_port, Q 
                           => n870);
   U2501 : NAND22 port map( A => n1362, B => position1_dp_cluster_7_N314, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_8_port);
   U2502 : NAND41 port map( A => position1_n868, B => position1_n869, C => 
                           position1_n870, D => position1_n871, Q => 
                           position1_n1589);
   U2503 : NAND22 port map( A => position1_y_sum_21_port, B => n511, Q => 
                           position1_n869);
   U2504 : NAND22 port map( A => position1_N1223_port, B => n639, Q => 
                           position1_n871);
   U2505 : AOI221 port map( A => position1_N556, B => n514, C => 
                           position1_N1000_port, D => n643, Q => position1_n870
                           );
   U2506 : NAND41 port map( A => position1_n864, B => position1_n865, C => 
                           position1_n866, D => position1_n867, Q => 
                           position1_n1588);
   U2507 : NAND22 port map( A => position1_y_sum_22_port, B => n511, Q => 
                           position1_n865);
   U2508 : NAND22 port map( A => position1_N1224_port, B => n639, Q => 
                           position1_n867);
   U2509 : AOI221 port map( A => position1_N557, B => n514, C => 
                           position1_N1001_port, D => n643, Q => position1_n866
                           );
   U2510 : NAND41 port map( A => position1_n972, B => position1_n973, C => 
                           position1_n974, D => position1_n975, Q => 
                           position1_n1615);
   U2511 : NAND22 port map( A => position1_x_sum_20_port, B => n510, Q => 
                           position1_n973);
   U2512 : NAND22 port map( A => position1_N1197_port, B => n637, Q => 
                           position1_n975);
   U2513 : AOI221 port map( A => position1_N505, B => n513, C => 
                           position1_N924_port, D => n641, Q => position1_n974)
                           ;
   U2514 : NAND41 port map( A => position1_n968, B => position1_n969, C => 
                           position1_n970, D => position1_n971, Q => 
                           position1_n1614);
   U2515 : NAND22 port map( A => position1_x_sum_21_port, B => n510, Q => 
                           position1_n969);
   U2516 : NAND22 port map( A => position1_N1198_port, B => n637, Q => 
                           position1_n971);
   U2517 : AOI221 port map( A => position1_N506, B => n513, C => 
                           position1_N925_port, D => n641, Q => position1_n970)
                           ;
   U2518 : INV3 port map( A => gensync1_n97, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port);
   U2519 : NAND22 port map( A => n816, B => gensync1_N139, Q => gensync1_n97);
   U2520 : XOR21 port map( A => gensync1_sub_91_2_cf_carry_2_port, B => 
                           gensync1_N171, Q => gensync1_N139);
   U2521 : NAND22 port map( A => gensync1_N174, B => n477, Q => gensync1_N85);
   U2522 : NOR21 port map( A => n396, B => n51, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_10_port);
   U2523 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_9_port,
                           Q => n396);
   U2524 : NOR21 port map( A => n381, B => n52, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_10_port);
   U2525 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_9_port,
                           Q => n381);
   U2526 : NOR21 port map( A => n398, B => n59, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_12_port);
   U2527 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_11_port
                           , Q => n398);
   U2528 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_5_port, Q 
                           => n862);
   U2529 : NAND22 port map( A => cam_x_5_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_5_port);
   U2530 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_1_port, Q 
                           => n809);
   U2531 : NOR21 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_0_port, B 
                           => n97, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_1_port);
   U2532 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_1_port);
   U2533 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_4_port, Q 
                           => n797);
   U2534 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_4_port);
   U2535 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_5_port, Q 
                           => n793);
   U2536 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_5_port);
   U2537 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_1_port, Q 
                           => n837);
   U2538 : NOR21 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_0_port, B 
                           => n98, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_1_port);
   U2539 : NAND22 port map( A => cam_x_1_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_1_port);
   U2540 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_1_port, Q 
                           => n836);
   U2541 : NOR21 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_0_port, B 
                           => n98, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_1_port);
   U2542 : NAND22 port map( A => cam_x_1_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_1_port);
   U2543 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_4_port, Q 
                           => n860);
   U2544 : NAND22 port map( A => cam_x_4_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_4_port);
   U2545 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_4_port, Q 
                           => n861);
   U2546 : NAND22 port map( A => cam_x_4_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_4_port);
   U2547 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_5_port, Q 
                           => n863);
   U2548 : NAND22 port map( A => cam_x_5_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_5_port);
   U2549 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_6_port, Q 
                           => n789);
   U2550 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_6_port);
   U2551 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_6_port, Q 
                           => n864);
   U2552 : NAND22 port map( A => cam_x_6_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_6_port);
   U2553 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_2_port, Q 
                           => n805);
   U2554 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_2_port);
   U2555 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_2_port, Q 
                           => n857);
   U2556 : NAND22 port map( A => n501, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_2_port);
   U2557 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_2_port, Q 
                           => n856);
   U2558 : NAND22 port map( A => cam_x_2_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_2_port);
   U2559 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_6_port, Q 
                           => n865);
   U2560 : NAND22 port map( A => cam_x_6_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_6_port);
   U2561 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_7_port, Q 
                           => n785);
   U2562 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_7_port);
   U2563 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_7_port, Q 
                           => n867);
   U2564 : NAND22 port map( A => cam_x_7_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_7_port);
   U2565 : INV3 port map( A => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_3_port, Q 
                           => n801);
   U2566 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => n1363, Q => 
                           position1_dp_cluster_5_mult_add_179_aco_PROD_not_3_port);
   U2567 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_3_port, Q 
                           => n859);
   U2568 : NAND22 port map( A => n499, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_3_port);
   U2569 : INV3 port map( A => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_3_port, Q 
                           => n858);
   U2570 : NAND22 port map( A => cam_x_3_port, B => n1363, Q => 
                           position1_dp_cluster_4_mult_add_178_aco_PROD_not_3_port);
   U2571 : INV3 port map( A => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_7_port, Q 
                           => n868);
   U2572 : NAND22 port map( A => cam_x_7_port, B => n1362, Q => 
                           position1_dp_cluster_0_mult_add_196_aco_PROD_not_7_port);
   U2573 : AOI221 port map( A => position1_N426, B => n646, C => position1_N653
                           , D => n649, Q => position1_n868);
   U2574 : XOR21 port map( A => position1_y_sum_21_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_21_port, Q 
                           => position1_N653);
   U2575 : XOR21 port map( A => position1_N376, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_21_port, Q 
                           => position1_N426);
   U2576 : AOI221 port map( A => position1_N427, B => n646, C => position1_N654
                           , D => n649, Q => position1_n864);
   U2577 : XOR21 port map( A => position1_y_sum_22_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_22_port, Q 
                           => position1_N654);
   U2578 : XOR21 port map( A => position1_N377, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_22_port, Q 
                           => position1_N427);
   U2579 : AOI221 port map( A => position1_N350_port, B => n644, C => 
                           position1_N627, D => n648, Q => position1_n972);
   U2580 : XOR21 port map( A => position1_x_sum_20_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_20_port, Q 
                           => position1_N627);
   U2581 : XOR21 port map( A => position1_N300, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_20_port, Q 
                           => position1_N350_port);
   U2582 : AOI221 port map( A => position1_N351_port, B => n644, C => 
                           position1_N628, D => n648, Q => position1_n968);
   U2583 : XOR21 port map( A => position1_x_sum_21_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_21_port, Q 
                           => position1_N628);
   U2584 : XOR21 port map( A => position1_N301, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_21_port, Q 
                           => position1_N351_port);
   U2585 : NOR21 port map( A => n507, B => n4, Q => n2134);
   U2586 : NOR21 port map( A => n507, B => n12, Q => n2133);
   U2587 : BUF2 port map( A => gensync1_N175, Q => n477);
   U2588 : NOR21 port map( A => n319, B => n52, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_10_port);
   U2589 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_9_port,
                           Q => n319);
   U2590 : NOR21 port map( A => n400, B => n58, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_14_port);
   U2591 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_13_port
                           , Q => n400);
   U2592 : NOR21 port map( A => n385, B => n65, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_14_port);
   U2593 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_13_port
                           , Q => n385);
   U2594 : NOR21 port map( A => n323, B => n65, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_14_port);
   U2595 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_13_port
                           , Q => n323);
   U2596 : NOR21 port map( A => n402, B => n57, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_16_port);
   U2597 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_15_port
                           , Q => n402);
   U2598 : NOR21 port map( A => n387, B => n64, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_16_port);
   U2599 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_15_port
                           , Q => n387);
   U2600 : NOR21 port map( A => n325, B => n64, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_16_port);
   U2601 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_15_port
                           , Q => n325);
   U2602 : NOR21 port map( A => n404, B => n56, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_18_port);
   U2603 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_17_port
                           , Q => n404);
   U2604 : NOR21 port map( A => n389, B => n63, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_18_port);
   U2605 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_17_port
                           , Q => n389);
   U2606 : NOR21 port map( A => n327, B => n63, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_18_port);
   U2607 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_17_port
                           , Q => n327);
   U2608 : NOR21 port map( A => n406, B => n55, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_20_port);
   U2609 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_19_port
                           , Q => n406);
   U2610 : NOR21 port map( A => n391, B => n62, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_20_port);
   U2611 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_19_port
                           , Q => n391);
   U2612 : NOR21 port map( A => n329, B => n62, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_20_port);
   U2613 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_19_port
                           , Q => n329);
   U2614 : NOR21 port map( A => n408, B => n54, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_22_port);
   U2615 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_21_port
                           , Q => n408);
   U2616 : NOR21 port map( A => n393, B => n61, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_22_port);
   U2617 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_21_port
                           , Q => n393);
   U2618 : NOR21 port map( A => n331, B => n61, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_22_port);
   U2619 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_21_port
                           , Q => n331);
   U2620 : XOR21 port map( A => position1_r409_carry_24_port, B => 
                           position1_y_sum_24_port, Q => position1_N379);
   U2621 : NOR21 port map( A => n210, B => n53, Q => 
                           position1_r409_carry_24_port);
   U2622 : INV3 port map( A => position1_r409_carry_23_port, Q => n210);
   U2623 : XOR21 port map( A => 
                           position1_dp_cluster_0_add_196_aco_carry_24_port, B 
                           => position1_x_sum_24_port, Q => 
                           position1_N1201_port);
   U2624 : NOR21 port map( A => n333, B => n60, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_24_port);
   U2625 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_23_port
                           , Q => n333);
   U2626 : NOR21 port map( A => n383, B => n66, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_12_port);
   U2627 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_11_port
                           , Q => n383);
   U2628 : NOR21 port map( A => n321, B => n66, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_12_port);
   U2629 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_11_port
                           , Q => n321);
   U2630 : NOR21 port map( A => n397, B => n69, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_11_port);
   U2631 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_10_port
                           , Q => n397);
   U2632 : NOR21 port map( A => n382, B => n70, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_11_port);
   U2633 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_10_port
                           , Q => n382);
   U2634 : NOR21 port map( A => n320, B => n70, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_11_port);
   U2635 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_10_port
                           , Q => n320);
   U2636 : NOR21 port map( A => n399, B => n76, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_13_port);
   U2637 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_12_port
                           , Q => n399);
   U2638 : NOR21 port map( A => n384, B => n82, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_13_port);
   U2639 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_12_port
                           , Q => n384);
   U2640 : NOR21 port map( A => n322, B => n82, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_13_port);
   U2641 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_12_port
                           , Q => n322);
   U2642 : NOR21 port map( A => n401, B => n75, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_15_port);
   U2643 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_14_port
                           , Q => n401);
   U2644 : NOR21 port map( A => n386, B => n81, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_15_port);
   U2645 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_14_port
                           , Q => n386);
   U2646 : NOR21 port map( A => n324, B => n81, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_15_port);
   U2647 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_14_port
                           , Q => n324);
   U2648 : NOR21 port map( A => n403, B => n74, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_17_port);
   U2649 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_16_port
                           , Q => n403);
   U2650 : NOR21 port map( A => n388, B => n80, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_17_port);
   U2651 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_16_port
                           , Q => n388);
   U2652 : NOR21 port map( A => n326, B => n80, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_17_port);
   U2653 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_16_port
                           , Q => n326);
   U2654 : NOR21 port map( A => n405, B => n73, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_19_port);
   U2655 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_18_port
                           , Q => n405);
   U2656 : NOR21 port map( A => n390, B => n79, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_19_port);
   U2657 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_18_port
                           , Q => n390);
   U2658 : NOR21 port map( A => n328, B => n79, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_19_port);
   U2659 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_18_port
                           , Q => n328);
   U2660 : NOR21 port map( A => n407, B => n72, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_21_port);
   U2661 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_20_port
                           , Q => n407);
   U2662 : NOR21 port map( A => n392, B => n78, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_21_port);
   U2663 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_20_port
                           , Q => n392);
   U2664 : NOR21 port map( A => n330, B => n78, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_21_port);
   U2665 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_20_port
                           , Q => n330);
   U2666 : NOR21 port map( A => n409, B => n71, Q => 
                           position1_dp_cluster_5_add_179_aco_carry_23_port);
   U2667 : INV3 port map( A => position1_dp_cluster_5_add_179_aco_carry_22_port
                           , Q => n409);
   U2668 : NOR21 port map( A => n394, B => n77, Q => 
                           position1_dp_cluster_4_add_178_aco_carry_23_port);
   U2669 : INV3 port map( A => position1_dp_cluster_4_add_178_aco_carry_22_port
                           , Q => n394);
   U2670 : NOR21 port map( A => n332, B => n77, Q => 
                           position1_dp_cluster_0_add_196_aco_carry_23_port);
   U2671 : INV3 port map( A => position1_dp_cluster_0_add_196_aco_carry_22_port
                           , Q => n332);
   U2672 : NAND31 port map( A => position1_n1147, B => position1_n357, C => 
                           position1_n1187, Q => position1_n1145);
   U2673 : NAND31 port map( A => position1_n1147, B => position1_gi_5_port, C 
                           => position1_n1187, Q => position1_n1151);
   U2674 : NOR40 port map( A => position1_n356, B => position1_n358, C => 
                           position1_gi_0_port, D => position1_gi_2_port, Q => 
                           position1_n1187);
   U2675 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_8_port, Q 
                           => n780);
   U2676 : NAND22 port map( A => n1362, B => position1_dp_cluster_6_N389, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_8_port);
   U2677 : NAND41 port map( A => position1_n880, B => position1_n881, C => 
                           position1_n882, D => position1_n883, Q => 
                           position1_n1592);
   U2678 : NAND22 port map( A => position1_y_sum_18_port, B => n511, Q => 
                           position1_n881);
   U2679 : NAND22 port map( A => position1_N1220_port, B => n639, Q => 
                           position1_n883);
   U2680 : AOI221 port map( A => position1_N553, B => n514, C => 
                           position1_N997_port, D => n643, Q => position1_n882)
                           ;
   U2681 : NAND41 port map( A => position1_n876, B => position1_n877, C => 
                           position1_n878, D => position1_n879, Q => 
                           position1_n1591);
   U2682 : NAND22 port map( A => position1_y_sum_19_port, B => n511, Q => 
                           position1_n877);
   U2683 : NAND22 port map( A => position1_N1221_port, B => n639, Q => 
                           position1_n879);
   U2684 : AOI221 port map( A => position1_N554, B => n514, C => 
                           position1_N998_port, D => n643, Q => position1_n878)
                           ;
   U2685 : NAND41 port map( A => position1_n872, B => position1_n873, C => 
                           position1_n874, D => position1_n875, Q => 
                           position1_n1590);
   U2686 : NAND22 port map( A => position1_y_sum_20_port, B => n511, Q => 
                           position1_n873);
   U2687 : NAND22 port map( A => position1_N1222_port, B => n639, Q => 
                           position1_n875);
   U2688 : AOI221 port map( A => position1_N555, B => n514, C => 
                           position1_N999_port, D => n643, Q => position1_n874)
                           ;
   U2689 : NAND41 port map( A => position1_n980, B => position1_n981, C => 
                           position1_n982, D => position1_n983, Q => 
                           position1_n1617);
   U2690 : NAND22 port map( A => position1_x_sum_18_port, B => n510, Q => 
                           position1_n981);
   U2691 : NAND22 port map( A => position1_N1195_port, B => n637, Q => 
                           position1_n983);
   U2692 : AOI221 port map( A => position1_N503, B => n513, C => 
                           position1_N922_port, D => n641, Q => position1_n982)
                           ;
   U2693 : NAND41 port map( A => position1_n976, B => position1_n977, C => 
                           position1_n978, D => position1_n979, Q => 
                           position1_n1616);
   U2694 : NAND22 port map( A => position1_x_sum_19_port, B => n510, Q => 
                           position1_n977);
   U2695 : NAND22 port map( A => position1_N1196_port, B => n637, Q => 
                           position1_n979);
   U2696 : AOI221 port map( A => position1_N504, B => n513, C => 
                           position1_N923_port, D => n641, Q => position1_n978)
                           ;
   U2697 : INV3 port map( A => gensync1_n96, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port);
   U2698 : NAND22 port map( A => n816, B => gensync1_N140, Q => gensync1_n96);
   U2699 : XOR21 port map( A => gensync1_sub_91_2_cf_carry_3_port, B => 
                           gensync1_N170, Q => gensync1_N140);
   U2700 : INV3 port map( A => gensync1_n95, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port);
   U2701 : NAND22 port map( A => n816, B => gensync1_N141, Q => gensync1_n95);
   U2702 : XOR21 port map( A => gensync1_sub_91_2_cf_carry_4_port, B => 
                           gensync1_N169, Q => gensync1_N141);
   U2703 : NOR21 port map( A => n336, B => n59, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_12_port);
   U2704 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_11_port
                           , Q => n336);
   U2705 : NOR21 port map( A => n9, B => n3, Q => 
                           gensync1_sub_91_2_cf_carry_2_port);
   U2706 : NOR21 port map( A => n8, B => n463, Q => 
                           gensync1_sub_91_2_cf_carry_3_port);
   U2707 : INV3 port map( A => gensync1_sub_91_2_cf_carry_2_port, Q => n463);
   U2708 : XOR21 port map( A => position1_y_sum_22_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_22_port, Q 
                           => position1_N1224_port);
   U2709 : XOR21 port map( A => position1_x_sum_22_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_22_port, Q 
                           => position1_N1199_port);
   U2710 : XOR21 port map( A => position1_y_sum_23_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_23_port, Q 
                           => position1_N1225_port);
   U2711 : XOR21 port map( A => position1_x_sum_23_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_23_port, Q 
                           => position1_N1200_port);
   U2712 : XOR21 port map( A => position1_x_sum_21_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_21_port, Q 
                           => position1_N1198_port);
   U2713 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_1_port, Q 
                           => n810);
   U2714 : NOR21 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_0_port, B 
                           => n97, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_1_port);
   U2715 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_1_port);
   U2716 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_4_port, Q 
                           => n798);
   U2717 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_5_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_4_port);
   U2718 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_5_port, Q 
                           => n794);
   U2719 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_6_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_5_port);
   U2720 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_2_port, Q 
                           => n806);
   U2721 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_3_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_2_port);
   U2722 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_6_port, Q 
                           => n790);
   U2723 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_6_port);
   U2724 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_3_port, Q 
                           => n802);
   U2725 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_3_port);
   U2726 : INV3 port map( A => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_7_port, Q 
                           => n786);
   U2727 : NAND22 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port, B 
                           => n1362, Q => 
                           position1_dp_cluster_1_mult_add_197_aco_PROD_not_7_port);
   U2728 : AOI221 port map( A => position1_N423, B => n646, C => position1_N650
                           , D => n649, Q => position1_n880);
   U2729 : XOR21 port map( A => position1_y_sum_18_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_18_port, Q 
                           => position1_N650);
   U2730 : XOR21 port map( A => position1_N373, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_18_port, Q 
                           => position1_N423);
   U2731 : AOI221 port map( A => position1_N424, B => n646, C => position1_N651
                           , D => n649, Q => position1_n876);
   U2732 : XOR21 port map( A => position1_y_sum_19_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_19_port, Q 
                           => position1_N651);
   U2733 : XOR21 port map( A => position1_N374, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_19_port, Q 
                           => position1_N424);
   U2734 : AOI221 port map( A => position1_N425, B => n646, C => position1_N652
                           , D => n649, Q => position1_n872);
   U2735 : XOR21 port map( A => position1_y_sum_20_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_20_port, Q 
                           => position1_N652);
   U2736 : XOR21 port map( A => position1_N375, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_20_port, Q 
                           => position1_N425);
   U2737 : AOI221 port map( A => position1_N348_port, B => n644, C => 
                           position1_N625, D => n648, Q => position1_n980);
   U2738 : XOR21 port map( A => position1_x_sum_18_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_18_port, Q 
                           => position1_N625);
   U2739 : XOR21 port map( A => position1_N298, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_18_port, Q 
                           => position1_N348_port);
   U2740 : AOI221 port map( A => position1_N349_port, B => n644, C => 
                           position1_N626, D => n648, Q => position1_n976);
   U2741 : XOR21 port map( A => position1_x_sum_19_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_19_port, Q 
                           => position1_N626);
   U2742 : XOR21 port map( A => position1_N299, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_19_port, Q 
                           => position1_N349_port);
   U2743 : NOR21 port map( A => n334, B => n51, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_10_port);
   U2744 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_9_port,
                           Q => n334);
   U2745 : NOR21 port map( A => n338, B => n58, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_14_port);
   U2746 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_13_port
                           , Q => n338);
   U2747 : NOR21 port map( A => n340, B => n57, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_16_port);
   U2748 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_15_port
                           , Q => n340);
   U2749 : NOR21 port map( A => n342, B => n56, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_18_port);
   U2750 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_17_port
                           , Q => n342);
   U2751 : NOR21 port map( A => n344, B => n55, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_20_port);
   U2752 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_19_port
                           , Q => n344);
   U2753 : NOR21 port map( A => n346, B => n54, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_22_port);
   U2754 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_21_port
                           , Q => n346);
   U2755 : XOR21 port map( A => 
                           position1_dp_cluster_1_add_197_aco_carry_24_port, B 
                           => position1_y_sum_24_port, Q => 
                           position1_N1226_port);
   U2756 : NOR21 port map( A => n348, B => n53, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_24_port);
   U2757 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_23_port
                           , Q => n348);
   U2758 : NOR21 port map( A => n335, B => n69, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_11_port);
   U2759 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_10_port
                           , Q => n335);
   U2760 : NOR21 port map( A => n337, B => n76, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_13_port);
   U2761 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_12_port
                           , Q => n337);
   U2762 : NOR21 port map( A => n339, B => n75, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_15_port);
   U2763 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_14_port
                           , Q => n339);
   U2764 : NOR21 port map( A => n341, B => n74, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_17_port);
   U2765 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_16_port
                           , Q => n341);
   U2766 : NOR21 port map( A => n343, B => n73, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_19_port);
   U2767 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_18_port
                           , Q => n343);
   U2768 : NOR21 port map( A => n345, B => n72, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_21_port);
   U2769 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_20_port
                           , Q => n345);
   U2770 : NOR21 port map( A => n347, B => n71, Q => 
                           position1_dp_cluster_1_add_197_aco_carry_23_port);
   U2771 : INV3 port map( A => position1_dp_cluster_1_add_197_aco_carry_22_port
                           , Q => n347);
   U2772 : NOR31 port map( A => position1_gi_3_port, B => position1_gi_7_port, 
                           C => position1_gi_1_port, Q => position1_n1147);
   U2773 : NAND41 port map( A => position1_n888, B => position1_n889, C => 
                           position1_n890, D => position1_n891, Q => 
                           position1_n1594);
   U2774 : NAND22 port map( A => position1_y_sum_16_port, B => n511, Q => 
                           position1_n889);
   U2775 : NAND22 port map( A => position1_N1218_port, B => n639, Q => 
                           position1_n891);
   U2776 : AOI221 port map( A => position1_N551, B => n514, C => 
                           position1_N995_port, D => n643, Q => position1_n890)
                           ;
   U2777 : NAND41 port map( A => position1_n884, B => position1_n885, C => 
                           position1_n886, D => position1_n887, Q => 
                           position1_n1593);
   U2778 : NAND22 port map( A => position1_y_sum_17_port, B => n511, Q => 
                           position1_n885);
   U2779 : NAND22 port map( A => position1_N1219_port, B => n639, Q => 
                           position1_n887);
   U2780 : AOI221 port map( A => position1_N552, B => n514, C => 
                           position1_N996_port, D => n643, Q => position1_n886)
                           ;
   U2781 : NAND41 port map( A => position1_n992, B => position1_n993, C => 
                           position1_n994, D => position1_n995, Q => 
                           position1_n1620);
   U2782 : NAND22 port map( A => position1_x_sum_15_port, B => n510, Q => 
                           position1_n993);
   U2783 : NAND22 port map( A => position1_N1192_port, B => n637, Q => 
                           position1_n995);
   U2784 : AOI221 port map( A => position1_N500, B => n513, C => 
                           position1_N919_port, D => n641, Q => position1_n994)
                           ;
   U2785 : NAND41 port map( A => position1_n988, B => position1_n989, C => 
                           position1_n990, D => position1_n991, Q => 
                           position1_n1619);
   U2786 : NAND22 port map( A => position1_x_sum_16_port, B => n510, Q => 
                           position1_n989);
   U2787 : NAND22 port map( A => position1_N1193_port, B => n637, Q => 
                           position1_n991);
   U2788 : AOI221 port map( A => position1_N501, B => n513, C => 
                           position1_N920_port, D => n641, Q => position1_n990)
                           ;
   U2789 : NAND41 port map( A => position1_n984, B => position1_n985, C => 
                           position1_n986, D => position1_n987, Q => 
                           position1_n1618);
   U2790 : NAND22 port map( A => position1_x_sum_17_port, B => n510, Q => 
                           position1_n985);
   U2791 : NAND22 port map( A => position1_N1194_port, B => n637, Q => 
                           position1_n987);
   U2792 : AOI221 port map( A => position1_N502, B => n513, C => 
                           position1_N921_port, D => n641, Q => position1_n986)
                           ;
   U2793 : INV3 port map( A => gensync1_n93, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_7_port);
   U2794 : NAND22 port map( A => n816, B => gensync1_N143, Q => gensync1_n93);
   U2795 : XNR21 port map( A => gensync1_sub_91_2_cf_carry_6_port, B => 
                           gensync1_N167, Q => gensync1_N143);
   U2796 : INV3 port map( A => gensync1_n92, Q => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_8_port);
   U2797 : NAND22 port map( A => n816, B => gensync1_N144, Q => gensync1_n92);
   U2798 : XNR21 port map( A => gensync1_sub_91_2_cf_carry_7_port, B => 
                           gensync1_N166, Q => gensync1_N144);
   U2799 : NAND22 port map( A => n816, B => gensync1_N142, Q => gensync1_n94);
   U2800 : XNR21 port map( A => gensync1_sub_91_2_cf_carry_5_port, B => 
                           gensync1_N168, Q => gensync1_N142);
   U2801 : NOR21 port map( A => n11, B => n464, Q => 
                           gensync1_sub_91_2_cf_carry_4_port);
   U2802 : INV3 port map( A => gensync1_sub_91_2_cf_carry_3_port, Q => n464);
   U2803 : XOR21 port map( A => position1_y_sum_20_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_20_port, Q 
                           => position1_N1222_port);
   U2804 : XOR21 port map( A => position1_x_sum_20_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_20_port, Q 
                           => position1_N1197_port);
   U2805 : XOR21 port map( A => position1_y_sum_21_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_21_port, Q 
                           => position1_N1223_port);
   U2806 : XOR21 port map( A => position1_x_sum_19_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_19_port, Q 
                           => position1_N1196_port);
   U2807 : AOI221 port map( A => position1_N421, B => n646, C => position1_N648
                           , D => n649, Q => position1_n888);
   U2808 : XOR21 port map( A => position1_y_sum_16_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_16_port, Q 
                           => position1_N648);
   U2809 : XOR21 port map( A => position1_N371, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_16_port, Q 
                           => position1_N421);
   U2810 : AOI221 port map( A => position1_N422, B => n646, C => position1_N649
                           , D => n649, Q => position1_n884);
   U2811 : XOR21 port map( A => position1_y_sum_17_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_17_port, Q 
                           => position1_N649);
   U2812 : XOR21 port map( A => position1_N372, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_17_port, Q 
                           => position1_N422);
   U2813 : AOI221 port map( A => position1_N345, B => n644, C => position1_N622
                           , D => n648, Q => position1_n992);
   U2814 : XOR21 port map( A => position1_x_sum_15_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_15_port, Q 
                           => position1_N622);
   U2815 : XOR21 port map( A => position1_N295, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_15_port, Q 
                           => position1_N345);
   U2816 : AOI221 port map( A => position1_N346_port, B => n644, C => 
                           position1_N623, D => n648, Q => position1_n988);
   U2817 : XOR21 port map( A => position1_x_sum_16_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_16_port, Q 
                           => position1_N623);
   U2818 : XOR21 port map( A => position1_N296, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_16_port, Q 
                           => position1_N346_port);
   U2819 : AOI221 port map( A => position1_N347_port, B => n644, C => 
                           position1_N624, D => n648, Q => position1_n984);
   U2820 : XOR21 port map( A => position1_x_sum_17_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_17_port, Q 
                           => position1_N624);
   U2821 : XOR21 port map( A => position1_N297, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_17_port, Q 
                           => position1_N347_port);
   U2822 : NOR21 port map( A => n507, B => n14, Q => n2131);
   U2823 : INV3 port map( A => n162, Q => gensync1_sub_91_2_cf_carry_6_port);
   U2824 : NOR21 port map( A => gensync1_N168, B => 
                           gensync1_sub_91_2_cf_carry_5_port, Q => n162);
   U2825 : INV3 port map( A => n163, Q => gensync1_sub_91_2_cf_carry_7_port);
   U2826 : NOR21 port map( A => gensync1_N167, B => 
                           gensync1_sub_91_2_cf_carry_6_port, Q => n163);
   U2827 : NOR21 port map( A => n13, B => n465, Q => 
                           gensync1_sub_91_2_cf_carry_5_port);
   U2828 : INV3 port map( A => gensync1_sub_91_2_cf_carry_4_port, Q => n465);
   U2829 : NAND41 port map( A => position1_n896, B => position1_n897, C => 
                           position1_n898, D => position1_n899, Q => 
                           position1_n1596);
   U2830 : NAND22 port map( A => position1_y_sum_14_port, B => n511, Q => 
                           position1_n897);
   U2831 : NAND22 port map( A => position1_N1216_port, B => n639, Q => 
                           position1_n899);
   U2832 : AOI221 port map( A => position1_N549, B => n514, C => 
                           position1_N993_port, D => n643, Q => position1_n898)
                           ;
   U2833 : NAND41 port map( A => position1_n892, B => position1_n893, C => 
                           position1_n894, D => position1_n895, Q => 
                           position1_n1595);
   U2834 : NAND22 port map( A => position1_y_sum_15_port, B => n511, Q => 
                           position1_n893);
   U2835 : NAND22 port map( A => position1_N1217_port, B => n639, Q => 
                           position1_n895);
   U2836 : AOI221 port map( A => position1_N550, B => n514, C => 
                           position1_N994_port, D => n643, Q => position1_n894)
                           ;
   U2837 : NAND41 port map( A => position1_n1000, B => position1_n1001, C => 
                           position1_n1002, D => position1_n1003, Q => 
                           position1_n1622);
   U2838 : NAND22 port map( A => position1_x_sum_13_port, B => n510, Q => 
                           position1_n1001);
   U2839 : NAND22 port map( A => position1_N1190_port, B => n637, Q => 
                           position1_n1003);
   U2840 : AOI221 port map( A => position1_N498, B => n513, C => 
                           position1_N917_port, D => n641, Q => position1_n1002
                           );
   U2841 : NAND41 port map( A => position1_n996, B => position1_n997, C => 
                           position1_n998, D => position1_n999, Q => 
                           position1_n1621);
   U2842 : NAND22 port map( A => position1_x_sum_14_port, B => n510, Q => 
                           position1_n997);
   U2843 : NAND22 port map( A => position1_N1191_port, B => n637, Q => 
                           position1_n999);
   U2844 : AOI221 port map( A => position1_N499, B => n513, C => 
                           position1_N918_port, D => n641, Q => position1_n998)
                           ;
   U2845 : NOR21 port map( A => gensync1_N166, B => 
                           gensync1_sub_91_2_cf_carry_7_port, Q => n164);
   U2846 : INV3 port map( A => gensync1_n91, Q => position1_dp_cluster_6_N389);
   U2847 : NAND22 port map( A => n816, B => gensync1_N145, Q => gensync1_n91);
   U2848 : XNR21 port map( A => gensync1_N165, B => 
                           gensync1_sub_91_2_cf_carry_8_port, Q => 
                           gensync1_N145);
   U2849 : INV3 port map( A => n164, Q => gensync1_sub_91_2_cf_carry_8_port);
   U2850 : XOR21 port map( A => position1_y_sum_18_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_18_port, Q 
                           => position1_N1220_port);
   U2851 : XOR21 port map( A => position1_x_sum_18_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_18_port, Q 
                           => position1_N1195_port);
   U2852 : XOR21 port map( A => position1_y_sum_19_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_19_port, Q 
                           => position1_N1221_port);
   U2853 : XOR21 port map( A => position1_x_sum_17_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_17_port, Q 
                           => position1_N1194_port);
   U2854 : AOI221 port map( A => position1_N419, B => n646, C => position1_N646
                           , D => n649, Q => position1_n896);
   U2855 : XOR21 port map( A => position1_y_sum_14_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_14_port, Q 
                           => position1_N646);
   U2856 : XOR21 port map( A => position1_N369_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_14_port, Q 
                           => position1_N419);
   U2857 : AOI221 port map( A => position1_N420, B => n646, C => position1_N647
                           , D => n649, Q => position1_n892);
   U2858 : XOR21 port map( A => position1_y_sum_15_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_15_port, Q 
                           => position1_N647);
   U2859 : XOR21 port map( A => position1_N370_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_15_port, Q 
                           => position1_N420);
   U2860 : AOI221 port map( A => position1_N343, B => n644, C => position1_N620
                           , D => n648, Q => position1_n1000);
   U2861 : XOR21 port map( A => position1_x_sum_13_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_13_port, Q 
                           => position1_N620);
   U2862 : XOR21 port map( A => position1_N293, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_13_port, Q 
                           => position1_N343);
   U2863 : AOI221 port map( A => position1_N344_port, B => n644, C => 
                           position1_N621, D => n648, Q => position1_n996);
   U2864 : XOR21 port map( A => position1_x_sum_14_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_14_port, Q 
                           => position1_N621);
   U2865 : XOR21 port map( A => position1_N294, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_14_port, Q 
                           => position1_N344_port);
   U2866 : NOR21 port map( A => n507, B => n15, Q => n2129);
   U2867 : NAND41 port map( A => position1_n904, B => position1_n905, C => 
                           position1_n906, D => position1_n907, Q => 
                           position1_n1598);
   U2868 : NAND22 port map( A => position1_y_sum_12_port, B => n511, Q => 
                           position1_n905);
   U2869 : NAND22 port map( A => position1_N1214_port, B => n639, Q => 
                           position1_n907);
   U2870 : AOI221 port map( A => position1_N547, B => n742, C => 
                           position1_N991_port, D => n642, Q => position1_n906)
                           ;
   U2871 : NAND41 port map( A => position1_n900, B => position1_n901, C => 
                           position1_n902, D => position1_n903, Q => 
                           position1_n1597);
   U2872 : NAND22 port map( A => position1_y_sum_13_port, B => n511, Q => 
                           position1_n901);
   U2873 : NAND22 port map( A => position1_N1215_port, B => n639, Q => 
                           position1_n903);
   U2874 : AOI221 port map( A => position1_N548, B => n742, C => 
                           position1_N992_port, D => n642, Q => position1_n902)
                           ;
   U2875 : NAND41 port map( A => position1_n1008, B => position1_n1009, C => 
                           position1_n1010, D => position1_n1011, Q => 
                           position1_n1624);
   U2876 : NAND22 port map( A => position1_x_sum_11_port, B => n512, Q => 
                           position1_n1009);
   U2877 : NAND22 port map( A => position1_N1188_port, B => n640, Q => 
                           position1_n1011);
   U2878 : AOI221 port map( A => position1_N496, B => n742, C => 
                           position1_N915_port, D => n642, Q => position1_n1010
                           );
   U2879 : NAND41 port map( A => position1_n1004, B => position1_n1005, C => 
                           position1_n1006, D => position1_n1007, Q => 
                           position1_n1623);
   U2880 : NAND22 port map( A => position1_x_sum_12_port, B => n510, Q => 
                           position1_n1005);
   U2881 : NAND22 port map( A => position1_N1189_port, B => n637, Q => 
                           position1_n1007);
   U2882 : AOI221 port map( A => position1_N497, B => n742, C => 
                           position1_N916_port, D => n641, Q => position1_n1006
                           );
   U2883 : XOR21 port map( A => position1_y_sum_16_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_16_port, Q 
                           => position1_N1218_port);
   U2884 : XOR21 port map( A => position1_x_sum_16_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_16_port, Q 
                           => position1_N1193_port);
   U2885 : XOR21 port map( A => position1_y_sum_17_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_17_port, Q 
                           => position1_N1219_port);
   U2886 : XOR21 port map( A => position1_x_sum_15_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_15_port, Q 
                           => position1_N1192_port);
   U2887 : AOI221 port map( A => position1_N417, B => n645, C => position1_N644
                           , D => n648, Q => position1_n904);
   U2888 : XOR21 port map( A => position1_y_sum_12_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_12_port, Q 
                           => position1_N644);
   U2889 : XOR21 port map( A => position1_N367_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_12_port, Q 
                           => position1_N417);
   U2890 : AOI221 port map( A => position1_N418, B => n645, C => position1_N645
                           , D => n649, Q => position1_n900);
   U2891 : XOR21 port map( A => position1_y_sum_13_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_13_port, Q 
                           => position1_N645);
   U2892 : XOR21 port map( A => position1_N368_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_13_port, Q 
                           => position1_N418);
   U2893 : AOI221 port map( A => position1_N341, B => n646, C => position1_N618
                           , D => n647, Q => position1_n1008);
   U2894 : XOR21 port map( A => position1_x_sum_11_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_11_port, Q 
                           => position1_N618);
   U2895 : XOR21 port map( A => position1_N291, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_11_port, Q 
                           => position1_N341);
   U2896 : AOI221 port map( A => position1_N342, B => position1_n858, C => 
                           position1_N619, D => n647, Q => position1_n1004);
   U2897 : XOR21 port map( A => position1_x_sum_12_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_12_port, Q 
                           => position1_N619);
   U2898 : XOR21 port map( A => position1_N292, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_12_port, Q 
                           => position1_N342);
   U2899 : NAND41 port map( A => position1_n912, B => position1_n913, C => 
                           position1_n914, D => position1_n915, Q => 
                           position1_n1600);
   U2900 : NAND22 port map( A => position1_y_sum_10_port, B => n675, Q => 
                           position1_n913);
   U2901 : NAND22 port map( A => position1_N1212_port, B => n638, Q => 
                           position1_n915);
   U2902 : AOI221 port map( A => position1_N415, B => n645, C => position1_N642
                           , D => n647, Q => position1_n912);
   U2903 : NAND41 port map( A => position1_n908, B => position1_n909, C => 
                           position1_n910, D => position1_n911, Q => 
                           position1_n1599);
   U2904 : NAND22 port map( A => position1_y_sum_11_port, B => n511, Q => 
                           position1_n909);
   U2905 : NAND22 port map( A => position1_N1213_port, B => n639, Q => 
                           position1_n911);
   U2906 : AOI221 port map( A => position1_N546, B => n742, C => 
                           position1_N990_port, D => n642, Q => position1_n910)
                           ;
   U2907 : NAND41 port map( A => position1_n1012, B => position1_n1013, C => 
                           position1_n1014, D => position1_n1015, Q => 
                           position1_n1625);
   U2908 : NAND22 port map( A => position1_x_sum_10_port, B => n512, Q => 
                           position1_n1013);
   U2909 : NAND22 port map( A => position1_N1187_port, B => n640, Q => 
                           position1_n1015);
   U2910 : AOI221 port map( A => position1_N495, B => n742, C => 
                           position1_N914_port, D => n643, Q => position1_n1014
                           );
   U2911 : NAND41 port map( A => position1_n916, B => position1_n917, C => 
                           position1_n918, D => position1_n919, Q => 
                           position1_n1601);
   U2912 : NAND22 port map( A => position1_y_sum_9_port, B => n675, Q => 
                           position1_n917);
   U2913 : NAND22 port map( A => position1_N1211_port, B => n638, Q => 
                           position1_n919);
   U2914 : AOI221 port map( A => position1_N544, B => n742, C => 
                           position1_N988_port, D => n642, Q => position1_n918)
                           ;
   U2915 : NAND41 port map( A => position1_n1020, B => position1_n1021, C => 
                           position1_n1022, D => position1_n1023, Q => 
                           position1_n1627);
   U2916 : NAND22 port map( A => position1_x_sum_8_port, B => n512, Q => 
                           position1_n1021);
   U2917 : NAND22 port map( A => position1_N1185_port, B => n640, Q => 
                           position1_n1023);
   U2918 : AOI221 port map( A => position1_N493, B => n742, C => 
                           position1_N912_port, D => position1_n857, Q => 
                           position1_n1022);
   U2919 : NAND41 port map( A => position1_n1016, B => position1_n1017, C => 
                           position1_n1018, D => position1_n1019, Q => 
                           position1_n1626);
   U2920 : NAND22 port map( A => position1_x_sum_9_port, B => n512, Q => 
                           position1_n1017);
   U2921 : NAND22 port map( A => position1_N1186_port, B => n640, Q => 
                           position1_n1019);
   U2922 : AOI221 port map( A => position1_N494, B => n742, C => 
                           position1_N913_port, D => position1_n857, Q => 
                           position1_n1018);
   U2923 : AOI221 port map( A => position1_N414, B => n645, C => position1_N641
                           , D => n648, Q => position1_n916);
   U2924 : XOR21 port map( A => position1_y_sum_9_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_9_port, Q 
                           => position1_N641);
   U2925 : AOI221 port map( A => position1_N339, B => position1_n858, C => 
                           position1_N616, D => n647, Q => position1_n1016);
   U2926 : XOR21 port map( A => position1_x_sum_9_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_9_port, Q 
                           => position1_N616);
   U2927 : AOI221 port map( A => position1_N340, B => position1_n858, C => 
                           position1_N617, D => n647, Q => position1_n1012);
   U2928 : XOR21 port map( A => position1_x_sum_10_port, B => 
                           position1_dp_cluster_4_add_178_aco_carry_10_port, Q 
                           => position1_N617);
   U2929 : XOR21 port map( A => position1_N290, B => 
                           position1_dp_cluster_7_add_0_root_add_170_3_carry_10_port, Q 
                           => position1_N340);
   U2930 : XOR21 port map( A => position1_y_sum_14_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_14_port, Q 
                           => position1_N1216_port);
   U2931 : XOR21 port map( A => position1_x_sum_12_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_12_port, Q 
                           => position1_N1189_port);
   U2932 : XOR21 port map( A => position1_x_sum_14_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_14_port, Q 
                           => position1_N1191_port);
   U2933 : XOR21 port map( A => position1_y_sum_13_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_13_port, Q 
                           => position1_N1215_port);
   U2934 : XOR21 port map( A => position1_y_sum_15_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_15_port, Q 
                           => position1_N1217_port);
   U2935 : XOR21 port map( A => position1_x_sum_13_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_13_port, Q 
                           => position1_N1190_port);
   U2936 : AOI221 port map( A => position1_N416, B => n645, C => position1_N643
                           , D => n649, Q => position1_n908);
   U2937 : XOR21 port map( A => position1_y_sum_11_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_11_port, Q 
                           => position1_N643);
   U2938 : XOR21 port map( A => position1_N366_port, B => 
                           position1_dp_cluster_6_add_0_root_add_171_3_carry_11_port, Q 
                           => position1_N416);
   U2939 : INV3 port map( A => position1_n1153, Q => n713);
   U2940 : AOI221 port map( A => position1_N224, B => n483, C => 
                           position1_count_img_19_port, D => n485, Q => 
                           position1_n1153);
   U2941 : XOR21 port map( A => position1_add_161_carry_19_port, B => 
                           position1_count_img_19_port, Q => position1_N224);
   U2942 : NAND41 port map( A => position1_n924, B => position1_n925, C => 
                           position1_n926, D => position1_n927, Q => 
                           position1_n1603);
   U2943 : NAND22 port map( A => position1_y_sum_7_port, B => n675, Q => 
                           position1_n925);
   U2944 : NAND22 port map( A => position1_N1209_port, B => n638, Q => 
                           position1_n927);
   U2945 : AOI221 port map( A => position1_N542, B => n742, C => 
                           position1_N986_port, D => n642, Q => position1_n926)
                           ;
   U2946 : NAND41 port map( A => position1_n920, B => position1_n921, C => 
                           position1_n922, D => position1_n923, Q => 
                           position1_n1602);
   U2947 : NAND22 port map( A => position1_y_sum_8_port, B => n675, Q => 
                           position1_n921);
   U2948 : NAND22 port map( A => position1_N1210_port, B => n638, Q => 
                           position1_n923);
   U2949 : AOI221 port map( A => position1_N543, B => n742, C => 
                           position1_N987_port, D => n642, Q => position1_n922)
                           ;
   U2950 : NAND41 port map( A => position1_n1024, B => position1_n1025, C => 
                           position1_n1026, D => position1_n1027, Q => 
                           position1_n1628);
   U2951 : NAND22 port map( A => position1_x_sum_7_port, B => n512, Q => 
                           position1_n1025);
   U2952 : NAND22 port map( A => position1_N1184_port, B => n640, Q => 
                           position1_n1027);
   U2953 : AOI221 port map( A => position1_N492, B => n742, C => 
                           position1_N911_port, D => position1_n857, Q => 
                           position1_n1026);
   U2954 : INV3 port map( A => position1_n1157, Q => n711);
   U2955 : AOI221 port map( A => position1_N222, B => position1_n1154, C => 
                           n484, D => position1_count_img_17_port, Q => 
                           position1_n1157);
   U2956 : XOR21 port map( A => position1_y_sum_12_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_12_port, Q 
                           => position1_N1214_port);
   U2957 : XOR21 port map( A => position1_x_sum_10_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_10_port, Q 
                           => position1_N1187_port);
   U2958 : XOR21 port map( A => position1_y_sum_11_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_11_port, Q 
                           => position1_N1213_port);
   U2959 : XOR21 port map( A => position1_x_sum_11_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_11_port, Q 
                           => position1_N1188_port);
   U2960 : XOR21 port map( A => position1_y_sum_10_port, B => 
                           position1_dp_cluster_5_add_179_aco_carry_10_port, Q 
                           => position1_N642);
   U2961 : BUF2 port map( A => position1_N560, Q => n516);
   U2962 : BUF2 port map( A => position1_N2460, Q => n633);
   U2963 : BUF2 port map( A => position1_N2459, Q => n629);
   U2964 : INV3 port map( A => position1_n1156, Q => n712);
   U2965 : AOI221 port map( A => position1_N223, B => n482, C => 
                           position1_count_img_18_port, D => n485, Q => 
                           position1_n1156);
   U2966 : NAND41 port map( A => position1_n928, B => position1_n929, C => 
                           position1_n930, D => position1_n931, Q => 
                           position1_n1604);
   U2967 : NAND22 port map( A => position1_y_sum_6_port, B => n675, Q => 
                           position1_n929);
   U2968 : NAND22 port map( A => position1_N1208_port, B => n638, Q => 
                           position1_n931);
   U2969 : AOI221 port map( A => position1_N541, B => n742, C => 
                           position1_N985_port, D => n642, Q => position1_n930)
                           ;
   U2970 : NAND41 port map( A => position1_n1032, B => position1_n1033, C => 
                           position1_n1034, D => position1_n1035, Q => 
                           position1_n1630);
   U2971 : NAND22 port map( A => position1_x_sum_5_port, B => n512, Q => 
                           position1_n1033);
   U2972 : NAND22 port map( A => position1_N1182_port, B => n640, Q => 
                           position1_n1035);
   U2973 : AOI221 port map( A => position1_N490, B => n742, C => 
                           position1_N909_port, D => position1_n857, Q => 
                           position1_n1034);
   U2974 : NAND41 port map( A => position1_n1028, B => position1_n1029, C => 
                           position1_n1030, D => position1_n1031, Q => 
                           position1_n1629);
   U2975 : NAND22 port map( A => position1_x_sum_6_port, B => n512, Q => 
                           position1_n1029);
   U2976 : NAND22 port map( A => position1_N1183_port, B => n640, Q => 
                           position1_n1031);
   U2977 : AOI221 port map( A => position1_N491, B => n742, C => 
                           position1_N910_port, D => position1_n857, Q => 
                           position1_n1030);
   U2978 : XOR21 port map( A => position1_y_sum_10_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_10_port, Q 
                           => position1_N1212_port);
   U2979 : XOR21 port map( A => position1_y_sum_9_port, B => 
                           position1_dp_cluster_1_add_197_aco_carry_9_port, Q 
                           => position1_N1211_port);
   U2980 : XOR21 port map( A => position1_x_sum_9_port, B => 
                           position1_dp_cluster_0_add_196_aco_carry_9_port, Q 
                           => position1_N1186_port);
   U2981 : BUF2 port map( A => position1_N2458, Q => n625);
   U2982 : INV3 port map( A => position1_n1158, Q => n710);
   U2983 : AOI221 port map( A => position1_N221, B => n483, C => n485, D => 
                           position1_count_img_16_port, Q => position1_n1158);
   U2984 : NOR31 port map( A => n2127, B => position1_count_img_19_port, C => 
                           position1_count_img_18_port, Q => position1_N267);
   U2985 : AOI211 port map( A => n499, B => position1_n1390, C => 
                           position1_n1391, Q => position1_n1389);
   U2986 : NOR31 port map( A => n2126, B => n2125, C => n18, Q => n2127);
   U2987 : NAND41 port map( A => position1_N2402, B => position1_N2391, C => 
                           position1_N2413, D => position1_n1579, Q => 
                           position1_n1182);
   U2988 : NAND41 port map( A => position1_n952, B => position1_n953, C => 
                           position1_n954, D => position1_n955, Q => 
                           position1_n1610);
   U2989 : NAND22 port map( A => position1_N1938, B => n675, Q => 
                           position1_n953);
   U2990 : AOI221 port map( A => position1_N355, B => n644, C => position1_N632
                           , D => n648, Q => position1_n952);
   U2991 : NAND22 port map( A => position1_N1202_port, B => n638, Q => 
                           position1_n955);
   U2992 : NAND41 port map( A => position1_n1052, B => position1_n1053, C => 
                           position1_n1054, D => position1_n1055, Q => 
                           position1_n1635);
   U2993 : NAND22 port map( A => position1_N1521_port, B => n512, Q => 
                           position1_n1053);
   U2994 : AOI221 port map( A => position1_N280, B => position1_n858, C => 
                           position1_N607, D => n647, Q => position1_n1052);
   U2995 : NAND22 port map( A => position1_N1177_port, B => n640, Q => 
                           position1_n1055);
   U2996 : NAND41 port map( A => position1_n948, B => position1_n949, C => 
                           position1_n950, D => position1_n951, Q => 
                           position1_n1609);
   U2997 : NAND22 port map( A => position1_y_sum_1_port, B => n675, Q => 
                           position1_n949);
   U2998 : AOI221 port map( A => position1_N406, B => n645, C => position1_N633
                           , D => position1_n859, Q => position1_n948);
   U2999 : NAND22 port map( A => position1_N1203_port, B => n638, Q => 
                           position1_n951);
   U3000 : NAND41 port map( A => position1_n1048, B => position1_n1049, C => 
                           position1_n1050, D => position1_n1051, Q => 
                           position1_n1634);
   U3001 : NAND22 port map( A => position1_x_sum_1_port, B => n512, Q => 
                           position1_n1049);
   U3002 : AOI221 port map( A => position1_N331, B => position1_n858, C => 
                           position1_N608, D => n647, Q => position1_n1048);
   U3003 : NAND22 port map( A => position1_N1178_port, B => n640, Q => 
                           position1_n1051);
   U3004 : NAND41 port map( A => position1_n944, B => position1_n945, C => 
                           position1_n946, D => position1_n947, Q => 
                           position1_n1608);
   U3005 : NAND22 port map( A => position1_y_sum_2_port, B => n675, Q => 
                           position1_n945);
   U3006 : AOI221 port map( A => position1_N407, B => n645, C => position1_N634
                           , D => position1_n859, Q => position1_n944);
   U3007 : NAND22 port map( A => position1_N1204_port, B => n638, Q => 
                           position1_n947);
   U3008 : NAND41 port map( A => position1_n940, B => position1_n941, C => 
                           position1_n942, D => position1_n943, Q => 
                           position1_n1607);
   U3009 : NAND22 port map( A => position1_y_sum_3_port, B => n675, Q => 
                           position1_n941);
   U3010 : AOI221 port map( A => position1_N408, B => n645, C => position1_N635
                           , D => position1_n859, Q => position1_n940);
   U3011 : NAND22 port map( A => position1_N1205_port, B => n638, Q => 
                           position1_n943);
   U3012 : NAND41 port map( A => position1_n936, B => position1_n937, C => 
                           position1_n938, D => position1_n939, Q => 
                           position1_n1606);
   U3013 : NAND22 port map( A => position1_y_sum_4_port, B => n675, Q => 
                           position1_n937);
   U3014 : AOI221 port map( A => position1_N409, B => n645, C => position1_N636
                           , D => position1_n859, Q => position1_n936);
   U3015 : NAND22 port map( A => position1_N1206_port, B => n638, Q => 
                           position1_n939);
   U3016 : NAND41 port map( A => position1_n932, B => position1_n933, C => 
                           position1_n934, D => position1_n935, Q => 
                           position1_n1605);
   U3017 : NAND22 port map( A => position1_y_sum_5_port, B => n675, Q => 
                           position1_n933);
   U3018 : NAND22 port map( A => position1_N1207_port, B => n638, Q => 
                           position1_n935);
   U3019 : AOI221 port map( A => position1_N410, B => n645, C => position1_N637
                           , D => position1_n859, Q => position1_n932);
   U3020 : NAND41 port map( A => position1_n1044, B => position1_n1045, C => 
                           position1_n1046, D => position1_n1047, Q => 
                           position1_n1633);
   U3021 : NAND22 port map( A => position1_x_sum_2_port, B => n512, Q => 
                           position1_n1045);
   U3022 : AOI221 port map( A => position1_N332, B => position1_n858, C => 
                           position1_N609, D => n647, Q => position1_n1044);
   U3023 : NAND22 port map( A => position1_N1179_port, B => n640, Q => 
                           position1_n1047);
   U3024 : NAND41 port map( A => position1_n1040, B => position1_n1041, C => 
                           position1_n1042, D => position1_n1043, Q => 
                           position1_n1632);
   U3025 : NAND22 port map( A => position1_x_sum_3_port, B => n675, Q => 
                           position1_n1041);
   U3026 : AOI221 port map( A => position1_N333, B => position1_n858, C => 
                           position1_N610, D => n647, Q => position1_n1040);
   U3027 : NAND22 port map( A => position1_N1180_port, B => n639, Q => 
                           position1_n1043);
   U3028 : NAND41 port map( A => position1_n1036, B => position1_n1037, C => 
                           position1_n1038, D => position1_n1039, Q => 
                           position1_n1631);
   U3029 : NAND22 port map( A => position1_x_sum_4_port, B => n675, Q => 
                           position1_n1037);
   U3030 : NAND22 port map( A => position1_N1181_port, B => n638, Q => 
                           position1_n1039);
   U3031 : AOI221 port map( A => position1_N334, B => n645, C => position1_N611
                           , D => n647, Q => position1_n1036);
   U3032 : INV3 port map( A => position1_n1160, Q => n708);
   U3033 : AOI221 port map( A => position1_N219, B => position1_n1154, C => 
                           position1_count_img_14_port, D => n484, Q => 
                           position1_n1160);
   U3034 : AOI221 port map( A => n1391, B => Y_barycentre_top_0_port, C => 
                           Y_barycentre_top_1_port, D => position1_N2383, Q => 
                           n1393);
   U3035 : AOI211 port map( A => position1_N2405, B => n23, C => gensync1_n99, 
                           Q => n1391);
   U3036 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_2_port, B 
                           => cam_y_0_port, Q => position1_N2405);
   U3037 : NOR21 port map( A => X_barycentre_top_6_port, B => n848, Q => n1446)
                           ;
   U3038 : INV3 port map( A => position1_N2378, Q => n848);
   U3039 : INV3 port map( A => position1_n1178, Q => n717);
   U3040 : AOI211 port map( A => reset_top, B => position1_gi_7_port, C => 
                           position1_n1179, Q => position1_n1178);
   U3041 : INV3 port map( A => position1_n1180, Q => n716);
   U3042 : AOI211 port map( A => reset_top, B => position1_gi_3_port, C => 
                           position1_n1179, Q => position1_n1180);
   U3043 : INV3 port map( A => position1_n1181, Q => n715);
   U3044 : AOI211 port map( A => reset_top, B => position1_gi_1_port, C => 
                           position1_n1179, Q => position1_n1181);
   U3045 : AOI2111 port map( A => position1_n1580, B => position1_n1581, C => 
                           n845, D => position1_n1582, Q => position1_n1579);
   U3046 : NOR40 port map( A => Y_barycentre_top_3_port, B => 
                           Y_barycentre_top_2_port, C => 
                           Y_barycentre_top_1_port, D => 
                           Y_barycentre_top_0_port, Q => position1_n1580);
   U3047 : NOR40 port map( A => Y_barycentre_top_6_port, B => n880, C => 
                           Y_barycentre_top_5_port, D => 
                           Y_barycentre_top_4_port, Q => position1_n1581);
   U3048 : NOR40 port map( A => n881, B => n882, C => X_barycentre_top_5_port, 
                           D => X_barycentre_top_4_port, Q => position1_n1582);
   U3049 : NOR21 port map( A => position1_n1177, B => position1_n368, Q => 
                           position1_N99);
   U3050 : NOR21 port map( A => position1_n1177, B => position1_n369, Q => 
                           position1_N98);
   U3051 : NOR21 port map( A => position1_n1177, B => position1_n370, Q => 
                           position1_N97);
   U3052 : NOR21 port map( A => position1_n1177, B => position1_n346, Q => 
                           position1_N88);
   U3053 : NOR21 port map( A => position1_n1177, B => position1_n347, Q => 
                           position1_N87);
   U3054 : NOR21 port map( A => position1_n1177, B => position1_n348, Q => 
                           position1_N86);
   U3055 : NOR21 port map( A => position1_n1177, B => position1_n349, Q => 
                           position1_N85);
   U3056 : NOR21 port map( A => position1_n1177, B => position1_n350, Q => 
                           position1_N84);
   U3057 : NOR21 port map( A => position1_n1177, B => position1_n351, Q => 
                           position1_N83);
   U3058 : NOR21 port map( A => position1_n1177, B => position1_n352, Q => 
                           position1_N82);
   U3059 : NOR21 port map( A => position1_n1177, B => position1_n353, Q => 
                           position1_N81);
   U3060 : NOR21 port map( A => position1_n1177, B => position1_n363, Q => 
                           position1_N104);
   U3061 : NOR21 port map( A => position1_n1177, B => position1_n364, Q => 
                           position1_N103);
   U3062 : NOR21 port map( A => position1_n1177, B => position1_n365, Q => 
                           position1_N102);
   U3063 : NOR21 port map( A => position1_n1177, B => position1_n366, Q => 
                           position1_N101);
   U3064 : NOR21 port map( A => position1_n1177, B => position1_n367, Q => 
                           position1_N100);
   U3065 : AOI221 port map( A => position1_N2395, B => n16, C => n1408, D => 
                           n1407, Q => n1409);
   U3066 : INV3 port map( A => position1_N2396, Q => n843);
   U3067 : AOI221 port map( A => Y_barycentre_top_2_port, B => n808, C => n1423
                           , D => n1422, Q => n1424);
   U3068 : NAND22 port map( A => position1_N2384, B => n21, Q => n1422);
   U3069 : INV3 port map( A => position1_N2384, Q => n808);
   U3070 : AOI221 port map( A => n1421, B => gensync1_n99, C => position1_N2383
                           , D => n23, Q => n1423);
   U3071 : AOI221 port map( A => X_barycentre_top_2_port, B => n852, C => n1438
                           , D => n1437, Q => n1439);
   U3072 : NAND22 port map( A => position1_N2374, B => n16, Q => n1437);
   U3073 : INV3 port map( A => position1_N2374, Q => n852);
   U3074 : INV3 port map( A => position1_N2385, Q => n804);
   U3075 : XNR21 port map( A => 
                           position1_dp_cluster_6_add_1_root_add_171_3_carry_4_port, B 
                           => position1_sub_250_3_carry_3_port, Q => 
                           position1_N2385);
   U3076 : AOI221 port map( A => n1436, B => n467, C => position1_N2373, D => 
                           n17, Q => n1438);
   U3077 : AOI211 port map( A => X_barycentre_top_1_port, B => position1_N2394,
                           C => X_barycentre_top_0_port, Q => n1436);
   U3078 : XOR21 port map( A => n503, B => cam_x_0_port, Q => position1_N2373);
   U3079 : NOR21 port map( A => Y_barycentre_top_7_port, B => n787, Q => n1403)
                           ;
   U3080 : NOR21 port map( A => position1_N2410, B => n31, Q => n1401);
   U3081 : AOI221 port map( A => n1406, B => X_barycentre_top_0_port, C => 
                           X_barycentre_top_1_port, D => position1_N2373, Q => 
                           n1408);
   U3082 : AOI211 port map( A => position1_N2394, B => n17, C => n467, Q => 
                           n1406);
   U3083 : XNR21 port map( A => n503, B => cam_x_0_port, Q => position1_N2394);
   U3084 : NOR21 port map( A => X_barycentre_top_5_port, B => n841, Q => n1414)
                           ;
   U3085 : NOR21 port map( A => position1_N2397, B => n20, Q => n1412);
   U3086 : NOR21 port map( A => Y_barycentre_top_5_port, B => n795, Q => n1399)
                           ;
   U3087 : NOR21 port map( A => position1_N2408, B => n26, Q => n1397);
   U3088 : NOR21 port map( A => X_barycentre_top_4_port, B => n850, Q => n1442)
                           ;
   U3089 : INV3 port map( A => position1_N2375, Q => n851);
   U3090 : NOR21 port map( A => Y_barycentre_top_4_port, B => n800, Q => n1427)
                           ;
   U3091 : INV3 port map( A => position1_N2386, Q => n800);
   U3092 : NOR21 port map( A => X_barycentre_top_7_port, B => n839, Q => n1418)
                           ;
   U3093 : NOR21 port map( A => position1_N2399, B => n25, Q => n1416);
   U3094 : BUF2 port map( A => position1_N2456, Q => n622);
   U3095 : INV3 port map( A => position1_N2387, Q => n796);
   U3096 : NOR21 port map( A => position1_N2387, B => n28, Q => n1429);
   U3097 : INV3 port map( A => position1_N2389, Q => n788);
   U3098 : NOR21 port map( A => position1_N2389, B => n32, Q => n1433);
   U3099 : NAND22 port map( A => Y_barycentre_top_2_port, B => n807, Q => n1392
                           );
   U3100 : INV3 port map( A => position1_N2406, Q => n807);
   U3101 : NOR21 port map( A => Y_barycentre_top_8_port, B => n782, Q => n1435)
                           ;
   U3102 : INV3 port map( A => position1_N2390, Q => n782);
   U3103 : NOR21 port map( A => Y_barycentre_top_6_port, B => n792, Q => n1431)
                           ;
   U3104 : INV3 port map( A => position1_N2388, Q => n792);
   U3105 : NAND22 port map( A => X_barycentre_top_2_port, B => n844, Q => n1407
                           );
   U3106 : INV3 port map( A => position1_N2395, Q => n844);
   U3107 : AOI221 port map( A => position1_N2406, B => n21, C => n1393, D => 
                           n1392, Q => n1394);
   U3108 : INV3 port map( A => position1_N2407, Q => n803);
   U3109 : INV3 port map( A => position1_N2381, Q => n845);
   U3110 : NOR21 port map( A => X_barycentre_top_8_port, B => n846, Q => n1450)
                           ;
   U3111 : AOI211 port map( A => Y_barycentre_top_1_port, B => position1_N2405,
                           C => Y_barycentre_top_0_port, Q => n1421);
   U3112 : INV3 port map( A => position1_n1159, Q => n709);
   U3113 : AOI221 port map( A => position1_N220, B => n482, C => n485, D => 
                           position1_count_img_15_port, Q => position1_n1159);
   U3114 : BUF2 port map( A => position1_N2460, Q => n632);
   U3115 : BUF2 port map( A => position1_N2455, Q => n470);
   U3116 : BUF2 port map( A => position1_N560, Q => n517);
   U3117 : BUF2 port map( A => position1_N2454, Q => n617);
   U3118 : INV3 port map( A => position1_n1162, Q => n706);
   U3119 : AOI221 port map( A => position1_N217, B => n482, C => 
                           position1_count_img_12_port, D => n485, Q => 
                           position1_n1162);
   U3120 : INV3 port map( A => position1_n1161, Q => n707);
   U3121 : AOI221 port map( A => position1_N218, B => n483, C => n485, D => 
                           position1_count_img_13_port, Q => position1_n1161);
   U3122 : INV3 port map( A => position1_n1163, Q => n705);
   U3123 : AOI221 port map( A => position1_N216, B => position1_n1154, C => 
                           n484, D => position1_count_img_11_port, Q => 
                           position1_n1163);
   U3124 : BUF2 port map( A => position1_N2458, Q => n623);
   U3125 : BUF2 port map( A => position1_N2459, Q => n627);
   U3126 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_7_port, C => image_process1_n89, Q
                           => image_process1_n86);
   U3127 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_3_port, C => image_process1_n89, Q
                           => image_process1_n106);
   U3128 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_1_port, C => image_process1_n89, Q
                           => image_process1_n114);
   U3129 : INV3 port map( A => image_process1_n88, Q => n774);
   U3130 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_7_port, C => image_process1_n89, Q
                           => image_process1_n88);
   U3131 : INV3 port map( A => image_process1_n108, Q => n770);
   U3132 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_3_port, C => image_process1_n89, Q
                           => image_process1_n108);
   U3133 : INV3 port map( A => image_process1_n116, Q => n768);
   U3134 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_1_port, C => image_process1_n89, Q
                           => image_process1_n116);
   U3135 : AOI211 port map( A => position1_count_img_13_port, B => n1355, C => 
                           position1_count_img_14_port, Q => n2125);
   U3136 : INV3 port map( A => n2124, Q => n1355);
   U3137 : AOI311 port map( A => position1_count_img_10_port, B => n1356, C => 
                           position1_count_img_11_port, D => 
                           position1_count_img_12_port, Q => n2124);
   U3138 : INV3 port map( A => n2123, Q => n1356);
   U3139 : AOI211 port map( A => position1_count_img_8_port, B => n2122, C => 
                           position1_count_img_9_port, Q => n2123);
   U3140 : NOR21 port map( A => position1_count_img_7_port, B => 
                           position1_count_img_6_port, Q => n2119);
   U3141 : NAND31 port map( A => position1_count_img_1_port, B => 
                           position1_count_img_0_port, C => 
                           position1_count_img_2_port, Q => n2121);
   U3142 : NAND31 port map( A => position1_count_img_4_port, B => 
                           position1_count_img_3_port, C => 
                           position1_count_img_5_port, Q => n2120);
   U3143 : XNR21 port map( A => gensync1_add_45_carry_9_port, B => 
                           gensync1_comptY_9_port, Q => n113);
   U3144 : BUF2 port map( A => position1_N2455, Q => n471);
   U3145 : BUF2 port map( A => position1_N2456, Q => n620);
   U3146 : BUF2 port map( A => position1_N2452, Q => n610);
   U3147 : NAND22 port map( A => image_process1_n86, B => image_process1_n87, Q
                           => image_process1_N31);
   U3148 : NAND22 port map( A => image_process1_bi_7_port, B => n490, Q => 
                           image_process1_n87);
   U3149 : NAND22 port map( A => image_process1_n106, B => image_process1_n107,
                           Q => image_process1_N19);
   U3150 : NAND22 port map( A => image_process1_bi_3_port, B => n490, Q => 
                           image_process1_n107);
   U3151 : NAND22 port map( A => image_process1_n114, B => image_process1_n115,
                           Q => image_process1_N13_port);
   U3152 : NAND22 port map( A => image_process1_bi_1_port, B => n490, Q => 
                           image_process1_n115);
   U3153 : NAND22 port map( A => image_process1_n86, B => image_process1_n90, Q
                           => image_process1_N29);
   U3154 : NAND22 port map( A => image_process1_ri_7_port, B => n490, Q => 
                           image_process1_n90);
   U3155 : NAND22 port map( A => image_process1_n106, B => image_process1_n109,
                           Q => image_process1_N17);
   U3156 : NAND22 port map( A => image_process1_ri_3_port, B => n490, Q => 
                           image_process1_n109);
   U3157 : NAND22 port map( A => image_process1_n114, B => image_process1_n118,
                           Q => image_process1_N11);
   U3158 : NAND22 port map( A => image_process1_ri_1_port, B => n490, Q => 
                           image_process1_n118);
   U3159 : INV3 port map( A => position1_n1165, Q => n703);
   U3160 : AOI221 port map( A => position1_N214, B => n482, C => 
                           position1_count_img_9_port, D => n485, Q => 
                           position1_n1165);
   U3161 : INV3 port map( A => position1_n1164, Q => n704);
   U3162 : AOI221 port map( A => position1_N215, B => n483, C => n485, D => 
                           position1_count_img_10_port, Q => position1_n1164);
   U3163 : NOR31 port map( A => image_process1_n27, B => SW1_top, C => 
                           gensync1_n103, Q => image_process1_n91);
   U3164 : AOI221 port map( A => image_process1_n56, B => image_process1_n57, C
                           => image_process1_gi_0_port, D => image_process1_n91
                           , Q => image_process1_n59);
   U3165 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_6_port, C => image_process1_n95, Q
                           => image_process1_n92);
   U3166 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_5_port, C => n778, Q => 
                           image_process1_n98);
   U3167 : AOI211 port map( A => image_process1_n91, B => 
                           image_process1_gi_4_port, C => n778, Q => 
                           image_process1_n102);
   U3168 : AOI221 port map( A => image_process1_n57, B => image_process1_n112, 
                           C => image_process1_n91, D => 
                           image_process1_gi_2_port, Q => image_process1_n110);
   U3169 : NOR21 port map( A => gensync1_n103, B => image_process1_state, Q => 
                           image_process1_n61);
   U3170 : INV3 port map( A => image_process1_n111, Q => n769);
   U3171 : AOI221 port map( A => image_process1_n57, B => image_process1_n112, 
                           C => image_process1_n58, D => 
                           image_process1_gi_2_port, Q => image_process1_n111);
   U3172 : XNR21 port map( A => gensync1_add_39_carry_9_port, B => 
                           gensync1_N174, Q => n114);
   U3173 : BUF2 port map( A => position1_N2452, Q => n609);
   U3174 : XOR21 port map( A => position1_N1938, B => n811, Q => position1_N632
                           );
   U3175 : XOR21 port map( A => position1_N1521_port, B => n854, Q => 
                           position1_N607);
   U3176 : BUF2 port map( A => position1_N2454, Q => n615);
   U3177 : BUF2 port map( A => position1_N2451, Q => n474);
   U3178 : BUF2 port map( A => position1_N2450, Q => n607);
   U3179 : NAND22 port map( A => image_process1_n92, B => image_process1_n93, Q
                           => image_process1_N28);
   U3180 : NAND22 port map( A => image_process1_bi_6_port, B => n490, Q => 
                           image_process1_n93);
   U3181 : NAND22 port map( A => image_process1_n98, B => image_process1_n99, Q
                           => image_process1_N25_port);
   U3182 : NAND22 port map( A => image_process1_bi_5_port, B => n490, Q => 
                           image_process1_n99);
   U3183 : NAND22 port map( A => image_process1_n102, B => image_process1_n103,
                           Q => image_process1_N22);
   U3184 : NAND22 port map( A => image_process1_bi_4_port, B => n490, Q => 
                           image_process1_n103);
   U3185 : NAND22 port map( A => image_process1_n92, B => image_process1_n96, Q
                           => image_process1_N26);
   U3186 : NAND22 port map( A => image_process1_ri_6_port, B => n490, Q => 
                           image_process1_n96);
   U3187 : NAND22 port map( A => image_process1_n98, B => image_process1_n101, 
                           Q => image_process1_N23);
   U3188 : NAND22 port map( A => image_process1_ri_5_port, B => n490, Q => 
                           image_process1_n101);
   U3189 : NAND22 port map( A => image_process1_n102, B => image_process1_n105,
                           Q => image_process1_N20);
   U3190 : NAND22 port map( A => image_process1_ri_4_port, B => n490, Q => 
                           image_process1_n105);
   U3191 : NAND22 port map( A => image_process1_n59, B => image_process1_n119, 
                           Q => image_process1_N10);
   U3192 : NAND22 port map( A => image_process1_bi_0_port, B => n490, Q => 
                           image_process1_n119);
   U3193 : NAND22 port map( A => image_process1_n59, B => image_process1_n60, Q
                           => image_process1_N8);
   U3194 : NAND22 port map( A => image_process1_ri_0_port, B => n490, Q => 
                           image_process1_n60);
   U3195 : INV3 port map( A => image_process1_n55, Q => n775);
   U3196 : AOI221 port map( A => image_process1_n56, B => image_process1_n57, C
                           => image_process1_n58, D => image_process1_gi_0_port
                           , Q => image_process1_n55);
   U3197 : INV3 port map( A => image_process1_n100, Q => n772);
   U3198 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_5_port, C => n778, Q => 
                           image_process1_n100);
   U3199 : INV3 port map( A => image_process1_n104, Q => n771);
   U3200 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_4_port, C => n778, Q => 
                           image_process1_n104);
   U3201 : INV3 port map( A => image_process1_n94, Q => n773);
   U3202 : AOI211 port map( A => image_process1_n58, B => 
                           image_process1_gi_6_port, C => image_process1_n95, Q
                           => image_process1_n94);
   U3203 : INV3 port map( A => position1_n1174, Q => n694);
   U3204 : AOI221 port map( A => position1_n802, B => n482, C => n485, D => 
                           position1_count_img_0_port, Q => position1_n1174);
   U3205 : INV3 port map( A => position1_n1173, Q => n695);
   U3206 : AOI221 port map( A => position1_N206, B => n483, C => n485, D => 
                           position1_count_img_1_port, Q => position1_n1173);
   U3207 : INV3 port map( A => position1_n1171, Q => n697);
   U3208 : AOI221 port map( A => position1_N208, B => n482, C => n484, D => 
                           position1_count_img_3_port, Q => position1_n1171);
   U3209 : INV3 port map( A => position1_n1170, Q => n698);
   U3210 : AOI221 port map( A => position1_N209, B => n483, C => n484, D => 
                           position1_count_img_4_port, Q => position1_n1170);
   U3211 : INV3 port map( A => position1_n1168, Q => n700);
   U3212 : AOI221 port map( A => position1_N211, B => n482, C => 
                           position1_count_img_6_port, D => n485, Q => 
                           position1_n1168);
   U3213 : INV3 port map( A => position1_n1167, Q => n701);
   U3214 : AOI221 port map( A => position1_N212, B => n483, C => 
                           position1_count_img_7_port, D => n485, Q => 
                           position1_n1167);
   U3215 : INV3 port map( A => position1_n1172, Q => n696);
   U3216 : AOI221 port map( A => position1_N207, B => position1_n1154, C => 
                           n485, D => position1_count_img_2_port, Q => 
                           position1_n1172);
   U3217 : INV3 port map( A => position1_n1169, Q => n699);
   U3218 : AOI221 port map( A => position1_N210, B => position1_n1154, C => 
                           n485, D => position1_count_img_5_port, Q => 
                           position1_n1169);
   U3219 : INV3 port map( A => position1_n1166, Q => n702);
   U3220 : AOI221 port map( A => position1_N213, B => position1_n1154, C => 
                           n485, D => position1_count_img_8_port, Q => 
                           position1_n1166);
   U3221 : NOR40 port map( A => position1_n1401, B => position1_n1402, C => 
                           n1354, D => n1352, Q => position1_n1144);
   U3222 : INV3 port map( A => position1_n1403, Q => n1352);
   U3223 : INV3 port map( A => position1_n1405, Q => n1354);
   U3224 : NAND41 port map( A => n1353, B => position1_count_img_16_port, C => 
                           position1_count_img_13_port, D => 
                           position1_count_img_15_port, Q => position1_n1402);
   U3225 : NAND41 port map( A => n1358, B => position1_count_img_4_port, C => 
                           position1_count_img_2_port, D => 
                           position1_count_img_3_port, Q => position1_n1401);
   U3226 : INV3 port map( A => position1_n1408, Q => n1358);
   U3227 : NAND22 port map( A => position1_count_img_8_port, B => 
                           position1_count_img_5_port, Q => position1_n1408);
   U3228 : NOR40 port map( A => position1_n1406, B => position1_n802, C => 
                           position1_count_img_14_port, D => 
                           position1_count_img_12_port, Q => position1_n1405);
   U3229 : NAND22 port map( A => position1_count_img_11_port, B => 
                           position1_count_img_10_port, Q => position1_n1406);
   U3230 : XOR21 port map( A => position1_N1938, B => n812, Q => 
                           position1_N1202_port);
   U3231 : XOR21 port map( A => position1_N1521_port, B => n855, Q => 
                           position1_N1177_port);
   U3232 : BUF2 port map( A => position1_N2451, Q => n473);
   U3233 : BUF2 port map( A => position1_N2450, Q => n606);
   U3234 : BUF2 port map( A => position1_N2448, Q => n603);
   U3235 : NOR40 port map( A => position1_count_img_6_port, B => n1357, C => 
                           position1_count_img_19_port, D => 
                           position1_count_img_18_port, Q => position1_n1403);
   U3236 : INV3 port map( A => position1_n1404, Q => n1357);
   U3237 : NOR21 port map( A => position1_count_img_7_port, B => 
                           position1_count_img_9_port, Q => position1_n1404);
   U3238 : NAND22 port map( A => position1_count_img_17_port, B => 
                           position1_count_img_16_port, Q => n2126);
   U3239 : INV3 port map( A => position1_n1407, Q => n1353);
   U3240 : NAND22 port map( A => position1_count_img_1_port, B => 
                           position1_count_img_17_port, Q => position1_n1407);
   U3241 : AOI2111 port map( A => image_process1_gi_5_port, B => n879, C => 
                           image_process1_gi_7_port, D => 
                           image_process1_gi_6_port, Q => 
                           image_process1_N62_port);
   U3242 : INV3 port map( A => n1388, Q => n879);
   U3243 : AOI2111 port map( A => image_process1_gi_2_port, B => 
                           image_process1_gi_1_port, C => 
                           image_process1_gi_4_port, D => 
                           image_process1_gi_3_port, Q => n1388);
   U3244 : NOR40 port map( A => position1_gi_2_port, B => position1_gi_4_port, 
                           C => position1_gi_5_port, D => position1_gi_6_port, 
                           Q => position1_n1148);
   U3245 : NAND31 port map( A => position1_n1147, B => position1_n362, C => 
                           position1_n1148, Q => position1_n1058);
   U3246 : AOI211 port map( A => image_process1_gi_6_port, B => n1387, C => 
                           image_process1_gi_7_port, Q => 
                           image_process1_N64_port);
   U3247 : NOR40 port map( A => image_process1_gi_3_port, B => 
                           image_process1_gi_2_port, C => 
                           image_process1_gi_1_port, D => 
                           image_process1_gi_0_port, Q => n1386);
   U3248 : NAND31 port map( A => position1_n1147, B => position1_gi_0_port, C 
                           => position1_n1148, Q => position1_n1065);
   U3249 : NOR40 port map( A => position1_n357, B => position1_n360, C => 
                           position1_n362, D => position1_gi_6_port, Q => 
                           position1_n1150);
   U3250 : NAND31 port map( A => position1_n1150, B => position1_n358, C => 
                           position1_n1147, Q => position1_n1146);
   U3251 : NAND31 port map( A => position1_n1147, B => position1_n1150, C => 
                           position1_gi_4_port, Q => position1_n1149);
   U3252 : NOR21 port map( A => position1_n344, B => position1_state_0_port, Q 
                           => position1_n1176);
   U3253 : BUF2 port map( A => position1_N2448, Q => n602);
   U3254 : NAND22 port map( A => position1_state_1_port, B => 
                           position1_state_0_port, Q => position1_n1152);
   U3255 : INV3 port map( A => reset_top, Q => n656);
   U3256 : NAND22 port map( A => n1389, B => n5, Q => n1390);
   U3257 : OAI311 port map( A => image_process1_gi_0_port, B => 
                           image_process1_gi_2_port, C => 
                           image_process1_gi_1_port, D => 
                           image_process1_gi_3_port, Q => n1389);
   U3258 : INV3 port map( A => position1_n1584, Q => n881);
   U3259 : NOR40 port map( A => X_barycentre_top_0_port, B => 
                           X_barycentre_top_1_port, C => 
                           X_barycentre_top_2_port, D => 
                           X_barycentre_top_3_port, Q => position1_n1584);
   U3260 : INV3 port map( A => position1_n1583, Q => n882);
   U3261 : NOR31 port map( A => X_barycentre_top_7_port, B => 
                           X_barycentre_top_8_port, C => 
                           X_barycentre_top_6_port, Q => position1_n1583);
   U3262 : NOR21 port map( A => n507, B => n34, Q => cam_x_9_port);
   U3263 : NOR31 port map( A => gensync1_N167, B => gensync1_N165, C => 
                           gensync1_N166, Q => n1374);
   U3264 : OAI311 port map( A => gensync1_N173, B => gensync1_N171, C => 
                           gensync1_N172, D => gensync1_N170, Q => n1375);
   U3265 : NOR31 port map( A => gensync1_N181, B => gensync1_N74, C => 
                           gensync1_N182, Q => gensync1_n90);
   U3266 : NAND22 port map( A => image_process1_state, B => SW1_top, Q => 
                           image_process1_n117);
   U3267 : NOR21 port map( A => n508, B => gensync1_N173, Q => gensync1_N56);
   U3268 : BUF2 port map( A => position1_N2445, Q => n594);
   U3269 : BUF2 port map( A => position1_N2446, Q => n598);
   U3270 : NOR41 port map( A => gensync1_n87, B => n875, C => n477, D => 
                           gensync1_N174, Q => gensync1_n107);
   U3271 : INV3 port map( A => gensync1_n88, Q => n875);
   U3272 : NAND22 port map( A => gensync1_n89, B => gensync1_n90, Q => 
                           gensync1_n87);
   U3273 : NOR31 port map( A => gensync1_N176, B => gensync1_N178, C => 
                           gensync1_N177, Q => gensync1_n88);
   U3274 : BUF2 port map( A => position1_N2446, Q => n599);
   U3275 : NAND22 port map( A => reset_top, B => gensync1_N43, Q => 
                           gensync1_n101);
   U3276 : NAND22 port map( A => gensync1_comptY_9_port, B => n1377, Q => 
                           gensync1_N43);
   U3277 : NAND31 port map( A => n1376, B => n1375, C => n1374, Q => n1377);
   U3278 : NOR21 port map( A => gensync1_N168, B => gensync1_N169, Q => n1376);
   U3279 : INV3 port map( A => reset_top, Q => n652);
   U3280 : BUF2 port map( A => position1_N2445, Q => n596);
   U3281 : INV3 port map( A => position1_n1585, Q => n880);
   U3282 : NOR21 port map( A => Y_barycentre_top_7_port, B => 
                           Y_barycentre_top_8_port, Q => position1_n1585);
   U3283 : INV3 port map( A => position1_N2353, Q => n1360);
   U3284 : INV3 port map( A => position1_n843, Q => n684);
   U3285 : AOI221 port map( A => n486, B => X_barycentre_top_8_port, C => n636,
                           D => position1_quot_x_8_port, Q => position1_n843);
   U3286 : INV3 port map( A => position1_n845, Q => n682);
   U3287 : AOI221 port map( A => n486, B => X_barycentre_top_6_port, C => n636,
                           D => position1_quot_x_6_port, Q => position1_n845);
   U3288 : INV3 port map( A => position1_n844, Q => n683);
   U3289 : AOI221 port map( A => n486, B => X_barycentre_top_7_port, C => n636,
                           D => position1_quot_x_7_port, Q => position1_n844);
   U3290 : INV3 port map( A => position1_n848, Q => n679);
   U3291 : AOI221 port map( A => n486, B => X_barycentre_top_3_port, C => n636,
                           D => position1_quot_x_3_port, Q => position1_n848);
   U3292 : INV3 port map( A => position1_n849, Q => n678);
   U3293 : AOI221 port map( A => n486, B => X_barycentre_top_2_port, C => n636,
                           D => position1_quot_x_2_port, Q => position1_n849);
   U3294 : INV3 port map( A => position1_n841, Q => n686);
   U3295 : AOI221 port map( A => n486, B => Y_barycentre_top_1_port, C => n636,
                           D => position1_quot_y_1_port, Q => position1_n841);
   U3296 : INV3 port map( A => position1_n850, Q => n677);
   U3297 : AOI221 port map( A => n486, B => X_barycentre_top_1_port, C => n636,
                           D => position1_quot_x_1_port, Q => position1_n850);
   U3298 : INV3 port map( A => position1_n842, Q => n685);
   U3299 : AOI221 port map( A => n486, B => Y_barycentre_top_0_port, C => n636,
                           D => position1_quot_y_0_port, Q => position1_n842);
   U3300 : INV3 port map( A => position1_n851, Q => n676);
   U3301 : AOI221 port map( A => n486, B => X_barycentre_top_0_port, C => n635,
                           D => position1_quot_x_0_port, Q => position1_n851);
   U3302 : AOI211 port map( A => n1359, B => position1_n1383, C => n654, Q => 
                           position1_N194);
   U3303 : NAND22 port map( A => position1_n344, B => position1_state_0_port, Q
                           => position1_n1383);
   U3304 : INV3 port map( A => position1_n1176, Q => n1359);
   U3305 : OAI2111 port map( A => gensync1_N178, B => n876, C => n477, D => 
                           gensync1_N174, Q => gensync1_N9);
   U3306 : INV3 port map( A => n1378, Q => n876);
   U3307 : NOR21 port map( A => gensync1_N176, B => gensync1_N177, Q => n1378);
   U3308 : INV3 port map( A => reset_top, Q => n655);
   U3309 : NOR21 port map( A => gensync1_N180, B => gensync1_N179, Q => 
                           gensync1_n89);
   U3310 : NOR21 port map( A => gensync1_n102, B => gensync1_N74, Q => 
                           gensync1_N22);
   U3311 : BUF2 port map( A => position1_N2452, Q => n612);
   U3312 : BUF2 port map( A => position1_N2460, Q => n631);
   U3313 : BUF2 port map( A => position1_N560, Q => n518);
   U3314 : INV3 port map( A => reset_top, Q => n654);
   U3315 : BUF2 port map( A => position1_N2446, Q => n600);
   U3316 : INV3 port map( A => reset_top, Q => n653);
   U3317 : BUF2 port map( A => position1_N2450, Q => n608);
   U3318 : BUF2 port map( A => position1_N2448, Q => n604);
   U3319 : BUF2 port map( A => position1_N2454, Q => n618);
   U3320 : INV3 port map( A => position1_n833, Q => n693);
   U3321 : AOI221 port map( A => n486, B => Y_barycentre_top_8_port, C => n636,
                           D => position1_quot_y_8_port, Q => position1_n833);
   U3322 : BUF2 port map( A => position1_N2460, Q => n634);
   U3323 : INV3 port map( A => position1_n847, Q => n680);
   U3324 : AOI221 port map( A => n486, B => X_barycentre_top_4_port, C => n635,
                           D => position1_quot_x_4_port, Q => position1_n847);
   U3325 : INV3 port map( A => position1_n838, Q => n689);
   U3326 : AOI221 port map( A => n486, B => Y_barycentre_top_4_port, C => n636,
                           D => position1_quot_y_4_port, Q => position1_n838);
   U3327 : INV3 port map( A => position1_n835, Q => n692);
   U3328 : AOI221 port map( A => n486, B => Y_barycentre_top_7_port, C => n636,
                           D => position1_quot_y_7_port, Q => position1_n835);
   U3329 : INV3 port map( A => position1_n836, Q => n691);
   U3330 : AOI221 port map( A => n486, B => Y_barycentre_top_6_port, C => n636,
                           D => position1_quot_y_6_port, Q => position1_n836);
   U3331 : INV3 port map( A => position1_n846, Q => n681);
   U3332 : AOI221 port map( A => n486, B => X_barycentre_top_5_port, C => 
                           position1_n834, D => position1_quot_x_5_port, Q => 
                           position1_n846);
   U3333 : INV3 port map( A => position1_n837, Q => n690);
   U3334 : AOI221 port map( A => n486, B => Y_barycentre_top_5_port, C => n636,
                           D => position1_quot_y_5_port, Q => position1_n837);
   U3335 : INV3 port map( A => position1_n839, Q => n688);
   U3336 : AOI221 port map( A => n486, B => Y_barycentre_top_3_port, C => n636,
                           D => position1_quot_y_3_port, Q => position1_n839);
   U3337 : INV3 port map( A => position1_n840, Q => n687);
   U3338 : AOI221 port map( A => n486, B => Y_barycentre_top_2_port, C => n636,
                           D => position1_quot_y_2_port, Q => position1_n840);
   U3339 : BUF2 port map( A => position1_N2456, Q => n621);
   U3340 : BUF2 port map( A => position1_N2459, Q => n628);
   U3341 : BUF2 port map( A => position1_N2445, Q => n595);
   U3342 : BUF2 port map( A => position1_N560, Q => n519);
   U3343 : INV3 port map( A => image_process1_n62, Q => n744);
   U3344 : NAND22 port map( A => reset_top, B => b_top(7), Q => 
                           image_process1_n62);
   U3345 : INV3 port map( A => position1_n1183, Q => n718);
   U3346 : NAND22 port map( A => b_out_proc_7_port, B => reset_top, Q => 
                           position1_n1183);
   U3347 : INV3 port map( A => position1_n1192, Q => n726);
   U3348 : NAND22 port map( A => g_out_proc_7_port, B => n651, Q => 
                           position1_n1192);
   U3349 : INV3 port map( A => position1_n1193, Q => n727);
   U3350 : NAND22 port map( A => g_out_proc_6_port, B => n651, Q => 
                           position1_n1193);
   U3351 : INV3 port map( A => position1_n1194, Q => n728);
   U3352 : NAND22 port map( A => g_out_proc_5_port, B => n651, Q => 
                           position1_n1194);
   U3353 : INV3 port map( A => position1_n1195, Q => n729);
   U3354 : NAND22 port map( A => g_out_proc_4_port, B => n651, Q => 
                           position1_n1195);
   U3355 : INV3 port map( A => position1_n1184, Q => n719);
   U3356 : NAND22 port map( A => b_out_proc_6_port, B => n651, Q => 
                           position1_n1184);
   U3357 : INV3 port map( A => position1_n1185, Q => n720);
   U3358 : NAND22 port map( A => b_out_proc_5_port, B => n651, Q => 
                           position1_n1185);
   U3359 : INV3 port map( A => position1_n1186, Q => n721);
   U3360 : NAND22 port map( A => b_out_proc_4_port, B => n651, Q => 
                           position1_n1186);
   U3361 : INV3 port map( A => position1_n1188, Q => n722);
   U3362 : NAND22 port map( A => b_out_proc_3_port, B => n651, Q => 
                           position1_n1188);
   U3363 : INV3 port map( A => position1_n1189, Q => n723);
   U3364 : NAND22 port map( A => b_out_proc_2_port, B => n651, Q => 
                           position1_n1189);
   U3365 : INV3 port map( A => position1_n1190, Q => n724);
   U3366 : NAND22 port map( A => b_out_proc_1_port, B => n651, Q => 
                           position1_n1190);
   U3367 : INV3 port map( A => position1_n1191, Q => n725);
   U3368 : NAND22 port map( A => b_out_proc_0_port, B => n651, Q => 
                           position1_n1191);
   U3369 : INV3 port map( A => position1_n1200, Q => n734);
   U3370 : NAND22 port map( A => r_out_proc_7_port, B => n651, Q => 
                           position1_n1200);
   U3371 : INV3 port map( A => position1_n1201, Q => n735);
   U3372 : NAND22 port map( A => r_out_proc_6_port, B => n651, Q => 
                           position1_n1201);
   U3373 : INV3 port map( A => position1_n1202, Q => n736);
   U3374 : NAND22 port map( A => r_out_proc_5_port, B => n651, Q => 
                           position1_n1202);
   U3375 : INV3 port map( A => position1_n1203, Q => n737);
   U3376 : NAND22 port map( A => r_out_proc_4_port, B => n651, Q => 
                           position1_n1203);
   U3377 : INV3 port map( A => position1_n1204, Q => n738);
   U3378 : NAND22 port map( A => r_out_proc_3_port, B => n651, Q => 
                           position1_n1204);
   U3379 : INV3 port map( A => position1_n1205, Q => n739);
   U3380 : NAND22 port map( A => r_out_proc_2_port, B => reset_top, Q => 
                           position1_n1205);
   U3381 : INV3 port map( A => position1_n1206, Q => n740);
   U3382 : NAND22 port map( A => r_out_proc_1_port, B => n651, Q => 
                           position1_n1206);
   U3383 : INV3 port map( A => position1_n1207, Q => n741);
   U3384 : NAND22 port map( A => r_out_proc_0_port, B => n651, Q => 
                           position1_n1207);
   U3385 : INV3 port map( A => position1_n1196, Q => n730);
   U3386 : NAND22 port map( A => g_out_proc_3_port, B => n651, Q => 
                           position1_n1196);
   U3387 : INV3 port map( A => position1_n1197, Q => n731);
   U3388 : NAND22 port map( A => g_out_proc_2_port, B => n651, Q => 
                           position1_n1197);
   U3389 : INV3 port map( A => position1_n1198, Q => n732);
   U3390 : NAND22 port map( A => g_out_proc_1_port, B => n651, Q => 
                           position1_n1198);
   U3391 : INV3 port map( A => position1_n1199, Q => n733);
   U3392 : NAND22 port map( A => g_out_proc_0_port, B => n651, Q => 
                           position1_n1199);
   U3393 : INV3 port map( A => image_process1_n70, Q => n752);
   U3394 : NAND22 port map( A => g_top(7), B => n650, Q => image_process1_n70);
   U3395 : INV3 port map( A => image_process1_n71, Q => n753);
   U3396 : NAND22 port map( A => g_top(6), B => n650, Q => image_process1_n71);
   U3397 : INV3 port map( A => image_process1_n72, Q => n754);
   U3398 : NAND22 port map( A => g_top(5), B => n650, Q => image_process1_n72);
   U3399 : INV3 port map( A => image_process1_n73, Q => n755);
   U3400 : NAND22 port map( A => g_top(4), B => n650, Q => image_process1_n73);
   U3401 : INV3 port map( A => image_process1_n63, Q => n745);
   U3402 : NAND22 port map( A => b_top(6), B => n650, Q => image_process1_n63);
   U3403 : INV3 port map( A => image_process1_n64, Q => n746);
   U3404 : NAND22 port map( A => b_top(5), B => n650, Q => image_process1_n64);
   U3405 : INV3 port map( A => image_process1_n65, Q => n747);
   U3406 : NAND22 port map( A => b_top(4), B => n650, Q => image_process1_n65);
   U3407 : INV3 port map( A => image_process1_n66, Q => n748);
   U3408 : NAND22 port map( A => b_top(3), B => n650, Q => image_process1_n66);
   U3409 : INV3 port map( A => image_process1_n67, Q => n749);
   U3410 : NAND22 port map( A => b_top(2), B => n650, Q => image_process1_n67);
   U3411 : INV3 port map( A => image_process1_n68, Q => n750);
   U3412 : NAND22 port map( A => b_top(1), B => n650, Q => image_process1_n68);
   U3413 : INV3 port map( A => image_process1_n69, Q => n751);
   U3414 : NAND22 port map( A => b_top(0), B => n650, Q => image_process1_n69);
   U3415 : INV3 port map( A => image_process1_n78, Q => n760);
   U3416 : NAND22 port map( A => r_top(7), B => reset_top, Q => 
                           image_process1_n78);
   U3417 : INV3 port map( A => image_process1_n79, Q => n761);
   U3418 : NAND22 port map( A => r_top(6), B => reset_top, Q => 
                           image_process1_n79);
   U3419 : INV3 port map( A => image_process1_n80, Q => n762);
   U3420 : NAND22 port map( A => r_top(5), B => reset_top, Q => 
                           image_process1_n80);
   U3421 : INV3 port map( A => image_process1_n81, Q => n763);
   U3422 : NAND22 port map( A => r_top(4), B => reset_top, Q => 
                           image_process1_n81);
   U3423 : INV3 port map( A => image_process1_n82, Q => n764);
   U3424 : NAND22 port map( A => r_top(3), B => reset_top, Q => 
                           image_process1_n82);
   U3425 : INV3 port map( A => image_process1_n83, Q => n765);
   U3426 : NAND22 port map( A => r_top(2), B => reset_top, Q => 
                           image_process1_n83);
   U3427 : INV3 port map( A => image_process1_n84, Q => n766);
   U3428 : NAND22 port map( A => r_top(1), B => reset_top, Q => 
                           image_process1_n84);
   U3429 : INV3 port map( A => image_process1_n85, Q => n767);
   U3430 : NAND22 port map( A => r_top(0), B => reset_top, Q => 
                           image_process1_n85);
   U3431 : INV3 port map( A => image_process1_n74, Q => n756);
   U3432 : NAND22 port map( A => g_top(3), B => reset_top, Q => 
                           image_process1_n74);
   U3433 : INV3 port map( A => image_process1_n75, Q => n757);
   U3434 : NAND22 port map( A => g_top(2), B => reset_top, Q => 
                           image_process1_n75);
   U3435 : INV3 port map( A => image_process1_n76, Q => n758);
   U3436 : NAND22 port map( A => g_top(1), B => reset_top, Q => 
                           image_process1_n76);
   U3437 : INV3 port map( A => image_process1_n77, Q => n759);
   U3438 : NAND22 port map( A => g_top(0), B => reset_top, Q => 
                           image_process1_n77);
   U3439 : NAND22 port map( A => position1_x_sum_7_port, B => n521, Q => 
                           position1_n1571);
   U3440 : NAND22 port map( A => position1_y_sum_7_port, B => n555, Q => 
                           position1_n1375);
   U3441 : NAND22 port map( A => position1_N1529_port, B => n521, Q => 
                           position1_n1570);
   U3442 : XNR21 port map( A => position1_x_sum_8_port, B => n515, Q => 
                           position1_N1529_port);
   U3443 : NAND22 port map( A => position1_N1946, B => n555, Q => 
                           position1_n1374);
   U3444 : XNR21 port map( A => position1_y_sum_8_port, B => n515, Q => 
                           position1_N1946);
   U3445 : NAND22 port map( A => position1_N1533_port, B => n521, Q => 
                           position1_n1566);
   U3446 : NAND22 port map( A => position1_N1950, B => n555, Q => 
                           position1_n1370);
   U3447 : NAND22 port map( A => position1_N1535_port, B => n520, Q => 
                           position1_n1564);
   U3448 : NAND22 port map( A => position1_N1952, B => n554, Q => 
                           position1_n1368);
   U3449 : NAND22 port map( A => position1_N1537_port, B => n520, Q => 
                           position1_n1562);
   U3450 : NAND22 port map( A => position1_N1954, B => n554, Q => 
                           position1_n1366);
   U3451 : NAND22 port map( A => position1_N1539_port, B => n520, Q => 
                           position1_n1560);
   U3452 : NAND22 port map( A => position1_N1956, B => n554, Q => 
                           position1_n1364);
   U3453 : NAND22 port map( A => position1_N1541_port, B => n520, Q => 
                           position1_n1558);
   U3454 : NAND22 port map( A => position1_N1958, B => n554, Q => 
                           position1_n1362);
   U3455 : NAND22 port map( A => position1_N1543_port, B => n520, Q => 
                           position1_n1556);
   U3456 : NAND22 port map( A => position1_N1960, B => n554, Q => 
                           position1_n1360);
   U3457 : NAND22 port map( A => position1_N1531_port, B => n521, Q => 
                           position1_n1568);
   U3458 : NAND22 port map( A => position1_N1948, B => n555, Q => 
                           position1_n1372);
   U3459 : NAND22 port map( A => position1_N1545_port, B => n520, Q => 
                           position1_n1554);
   U3460 : NAND22 port map( A => position1_N1962, B => n554, Q => 
                           position1_n1358);
   U3461 : AOI221 port map( A => position1_x_sum_12_port, B => n248, C => n2093
                           , D => n1342, Q => n2095);
   U3462 : INV3 port map( A => n2092, Q => n1342);
   U3463 : AOI221 port map( A => n2091, B => n1344, C => n625, D => n66, Q => 
                           n2093);
   U3464 : NOR21 port map( A => n276, B => position1_x_sum_12_port, Q => n2092)
                           ;
   U3465 : AOI221 port map( A => position1_y_sum_12_port, B => n42, C => n1759,
                           D => n1341, Q => n1761);
   U3466 : INV3 port map( A => n1758, Q => n1341);
   U3467 : AOI221 port map( A => n1757, B => n1343, C => n625, D => n59, Q => 
                           n1759);
   U3468 : NOR21 port map( A => n276, B => position1_y_sum_12_port, Q => n1758)
                           ;
   U3469 : AOI221 port map( A => position1_x_sum_14_port, B => n252, C => n2097
                           , D => n1338, Q => n2099);
   U3470 : INV3 port map( A => n2096, Q => n1338);
   U3471 : AOI221 port map( A => n2095, B => n1340, C => n622, D => n65, Q => 
                           n2097);
   U3472 : NOR21 port map( A => n46, B => position1_x_sum_14_port, Q => n2096);
   U3473 : AOI221 port map( A => position1_y_sum_14_port, B => n280, C => n1763
                           , D => n1337, Q => n1765);
   U3474 : INV3 port map( A => n1762, Q => n1337);
   U3475 : AOI221 port map( A => n1761, B => n1339, C => n622, D => n58, Q => 
                           n1763);
   U3476 : NOR21 port map( A => n280, B => position1_y_sum_14_port, Q => n1762)
                           ;
   U3477 : AOI221 port map( A => position1_x_sum_16_port, B => n284, C => n2101
                           , D => n1334, Q => n2103);
   U3478 : INV3 port map( A => n2100, Q => n1334);
   U3479 : AOI221 port map( A => n2099, B => n1336, C => n618, D => n64, Q => 
                           n2101);
   U3480 : NOR21 port map( A => n284, B => position1_x_sum_16_port, Q => n2100)
                           ;
   U3481 : AOI221 port map( A => position1_y_sum_16_port, B => n256, C => n1767
                           , D => n1333, Q => n1769);
   U3482 : INV3 port map( A => n1766, Q => n1333);
   U3483 : AOI221 port map( A => n1765, B => n1335, C => n618, D => n57, Q => 
                           n1767);
   U3484 : NOR21 port map( A => n256, B => position1_y_sum_16_port, Q => n1766)
                           ;
   U3485 : AOI221 port map( A => position1_x_sum_18_port, B => n288, C => n2105
                           , D => n1330, Q => n2107);
   U3486 : INV3 port map( A => n2104, Q => n1330);
   U3487 : AOI221 port map( A => n2103, B => n1332, C => n613, D => n63, Q => 
                           n2105);
   U3488 : NOR21 port map( A => n47, B => position1_x_sum_18_port, Q => n2104);
   U3489 : AOI221 port map( A => position1_y_sum_18_port, B => n259, C => n1771
                           , D => n1329, Q => n1773);
   U3490 : INV3 port map( A => n1770, Q => n1329);
   U3491 : AOI221 port map( A => n1769, B => n1331, C => n612, D => n56, Q => 
                           n1771);
   U3492 : NOR21 port map( A => n47, B => position1_y_sum_18_port, Q => n1770);
   U3493 : AOI221 port map( A => position1_x_sum_20_port, B => n263, C => n2109
                           , D => n1326, Q => n2111);
   U3494 : INV3 port map( A => n2108, Q => n1326);
   U3495 : AOI221 port map( A => n2107, B => n1328, C => n608, D => n62, Q => 
                           n2109);
   U3496 : NOR21 port map( A => n44, B => position1_x_sum_20_port, Q => n2108);
   U3497 : AOI221 port map( A => position1_y_sum_20_port, B => n292, C => n1775
                           , D => n1325, Q => n1777);
   U3498 : INV3 port map( A => n1774, Q => n1325);
   U3499 : AOI221 port map( A => n1773, B => n1327, C => n608, D => n55, Q => 
                           n1775);
   U3500 : NOR21 port map( A => n263, B => position1_y_sum_20_port, Q => n1774)
                           ;
   U3501 : AOI221 port map( A => position1_x_sum_22_port, B => n267, C => n2113
                           , D => n1322, Q => n2115);
   U3502 : INV3 port map( A => n2112, Q => n1322);
   U3503 : AOI221 port map( A => n2111, B => n1324, C => n604, D => n61, Q => 
                           n2113);
   U3504 : NOR21 port map( A => n43, B => position1_x_sum_22_port, Q => n2112);
   U3505 : AOI221 port map( A => position1_y_sum_22_port, B => n267, C => n1779
                           , D => n1321, Q => n1781);
   U3506 : INV3 port map( A => n1778, Q => n1321);
   U3507 : AOI221 port map( A => n1777, B => n1323, C => n604, D => n54, Q => 
                           n1779);
   U3508 : NOR21 port map( A => n296, B => position1_y_sum_22_port, Q => n1778)
                           ;
   U3509 : AOI221 port map( A => position1_x_sum_10_port, B => n272, C => n1346
                           , D => n2089, Q => n2091);
   U3510 : INV3 port map( A => n2088, Q => n1346);
   U3511 : NAND22 port map( A => n632, B => n52, Q => n2089);
   U3512 : AOI221 port map( A => position1_y_sum_10_port, B => n245, C => n1345
                           , D => n1755, Q => n1757);
   U3513 : INV3 port map( A => n1754, Q => n1345);
   U3514 : NAND22 port map( A => n633, B => n51, Q => n1755);
   U3515 : NOR40 port map( A => position1_x_sum_7_port, B => 
                           position1_x_sum_6_port, C => position1_x_sum_5_port,
                           D => position1_x_sum_4_port, Q => n2083);
   U3516 : NOR40 port map( A => position1_y_sum_7_port, B => 
                           position1_y_sum_6_port, C => position1_y_sum_5_port,
                           D => position1_y_sum_4_port, Q => n1749);
   U3517 : NAND22 port map( A => position1_x_sum_4_port, B => n521, Q => 
                           position1_n1574);
   U3518 : NAND22 port map( A => position1_y_sum_4_port, B => n555, Q => 
                           position1_n1378);
   U3519 : NAND22 port map( A => position1_x_sum_3_port, B => n521, Q => 
                           position1_n1575);
   U3520 : NAND22 port map( A => position1_y_sum_3_port, B => n555, Q => 
                           position1_n1379);
   U3521 : NAND22 port map( A => position1_x_sum_5_port, B => n521, Q => 
                           position1_n1573);
   U3522 : NAND22 port map( A => position1_y_sum_5_port, B => n555, Q => 
                           position1_n1377);
   U3523 : NAND22 port map( A => position1_x_sum_6_port, B => n521, Q => 
                           position1_n1572);
   U3524 : NAND22 port map( A => position1_y_sum_6_port, B => n555, Q => 
                           position1_n1376);
   U3525 : NAND22 port map( A => position1_N1521_port, B => n521, Q => 
                           position1_n1578);
   U3526 : NAND22 port map( A => position1_N1938, B => n555, Q => 
                           position1_n1382);
   U3527 : NAND22 port map( A => position1_x_sum_1_port, B => n522, Q => 
                           position1_n1577);
   U3528 : NAND22 port map( A => position1_y_sum_1_port, B => n556, Q => 
                           position1_n1381);
   U3529 : NAND22 port map( A => position1_x_sum_2_port, B => n521, Q => 
                           position1_n1576);
   U3530 : NAND22 port map( A => position1_y_sum_2_port, B => n555, Q => 
                           position1_n1380);
   U3531 : NOR21 port map( A => n588, B => n2118, Q => position1_N1519_port);
   U3532 : AOI221 port map( A => position1_x_sum_24_port, B => n300, C => n2117
                           , D => n1348, Q => n2118);
   U3533 : INV3 port map( A => n2116, Q => n1348);
   U3534 : AOI221 port map( A => n2115, B => n1320, C => n600, D => n60, Q => 
                           n2117);
   U3535 : NOR21 port map( A => n588, B => n1784, Q => position1_N1936);
   U3536 : AOI221 port map( A => position1_y_sum_24_port, B => n300, C => n1783
                           , D => n1347, Q => n1784);
   U3537 : INV3 port map( A => n1782, Q => n1347);
   U3538 : AOI221 port map( A => n1781, B => n1101, C => n600, D => n53, Q => 
                           n1783);
   U3539 : NOR21 port map( A => n300, B => position1_x_sum_24_port, Q => n2116)
                           ;
   U3540 : NOR21 port map( A => n300, B => position1_y_sum_24_port, Q => n1782)
                           ;
   U3541 : INV3 port map( A => n2085, Q => n1350);
   U3542 : AOI221 port map( A => n2084, B => n2083, C => n518, D => n50, Q => 
                           n2085);
   U3543 : NOR40 port map( A => position1_x_sum_3_port, B => 
                           position1_x_sum_2_port, C => position1_x_sum_1_port,
                           D => position1_N1521_port, Q => n2084);
   U3544 : INV3 port map( A => n1751, Q => n1349);
   U3545 : AOI221 port map( A => n1750, B => n1749, C => n518, D => n49, Q => 
                           n1751);
   U3546 : NOR40 port map( A => position1_y_sum_3_port, B => 
                           position1_y_sum_2_port, C => position1_y_sum_1_port,
                           D => position1_N1938, Q => n1750);
   U3547 : INV3 port map( A => n166, Q => position1_sub_216_carry_9_port);
   U3548 : NOR21 port map( A => n515, B => position1_x_sum_8_port, Q => n166);
   U3549 : INV3 port map( A => n165, Q => position1_sub_226_carry_9_port);
   U3550 : NOR21 port map( A => n515, B => position1_y_sum_8_port, Q => n165);
   U3551 : BUF2 port map( A => position1_N2452, Q => n611);
   U3552 : BUF2 port map( A => position1_N2445, Q => n593);
   U3553 : BUF2 port map( A => position1_N2459, Q => n626);
   U3554 : BUF2 port map( A => position1_N2456, Q => n619);
   U3555 : BUF2 port map( A => position1_N2450, Q => n605);
   U3556 : BUF2 port map( A => position1_N2448, Q => n601);
   U3557 : BUF2 port map( A => position1_N2458, Q => n624);
   U3558 : BUF2 port map( A => position1_N2446, Q => n597);
   U3559 : BUF2 port map( A => position1_N2454, Q => n614);
   U3560 : BUF2 port map( A => position1_N2454, Q => n616);
   U3561 : BUF2 port map( A => position1_N2452, Q => n613);
   U3562 : LOGIC1 port map( Q => position1_n283);
   U3563 : OAI212 port map( A => n1370, B => n1369, C => n1368, Q => n1371);
   U3564 : OAI212 port map( A => gensync1_N181, B => gensync1_N182, C => 
                           gensync1_N180, Q => n1380);
   U3565 : OAI212 port map( A => gensync1_N181, B => gensync1_N182, C => 
                           gensync1_N180, Q => n1382);
   U3566 : OAI212 port map( A => n1386, B => n5, C => n33, Q => n1387);
   U3567 : OAI212 port map( A => Y_barycentre_top_3_port, B => n803, C => n1394
                           , Q => n1395);
   U3568 : OAI212 port map( A => position1_N2407, B => n24, C => n1395, Q => 
                           n1396);
   U3569 : OAI222 port map( A => n1397, B => n1396, C => 
                           Y_barycentre_top_4_port, D => n799, Q => n1398);
   U3570 : OAI222 port map( A => position1_N2409, B => n28, C => n1399, D => 
                           n1398, Q => n1400);
   U3571 : OAI222 port map( A => n1401, B => n1400, C => 
                           Y_barycentre_top_6_port, D => n791, Q => n1402);
   U3572 : OAI222 port map( A => position1_N2411, B => n32, C => n1403, D => 
                           n1402, Q => n1404);
   U3573 : OAI222 port map( A => n1405, B => n1404, C => 
                           Y_barycentre_top_8_port, D => n781, Q => 
                           position1_N2413);
   U3574 : OAI212 port map( A => X_barycentre_top_3_port, B => n843, C => n1409
                           , Q => n1410);
   U3575 : OAI212 port map( A => position1_N2396, B => n19, C => n1410, Q => 
                           n1411);
   U3576 : OAI222 port map( A => n1412, B => n1411, C => 
                           X_barycentre_top_4_port, D => n842, Q => n1413);
   U3577 : OAI222 port map( A => position1_N2398, B => n22, C => n1414, D => 
                           n1413, Q => n1415);
   U3578 : OAI222 port map( A => n1416, B => n1415, C => 
                           X_barycentre_top_6_port, D => n840, Q => n1417);
   U3579 : OAI222 port map( A => position1_N2400, B => n27, C => n1418, D => 
                           n1417, Q => n1419);
   U3580 : OAI222 port map( A => n1420, B => n1419, C => 
                           X_barycentre_top_8_port, D => n838, Q => 
                           position1_N2402);
   U3581 : OAI212 port map( A => position1_N2385, B => n24, C => n1424, Q => 
                           n1425);
   U3582 : OAI212 port map( A => Y_barycentre_top_3_port, B => n804, C => n1425
                           , Q => n1426);
   U3583 : OAI222 port map( A => n1427, B => n1426, C => position1_N2386, D => 
                           n26, Q => n1428);
   U3584 : OAI222 port map( A => Y_barycentre_top_5_port, B => n796, C => n1429
                           , D => n1428, Q => n1430);
   U3585 : OAI222 port map( A => n1431, B => n1430, C => position1_N2388, D => 
                           n31, Q => n1432);
   U3586 : OAI222 port map( A => Y_barycentre_top_7_port, B => n788, C => n1433
                           , D => n1432, Q => n1434);
   U3587 : OAI222 port map( A => n1435, B => n1434, C => position1_N2390, D => 
                           n30, Q => position1_N2391);
   U3588 : OAI212 port map( A => position1_N2375, B => n19, C => n1439, Q => 
                           n1440);
   U3589 : OAI212 port map( A => X_barycentre_top_3_port, B => n851, C => n1440
                           , Q => n1441);
   U3590 : OAI222 port map( A => n1442, B => n1441, C => position1_N2376, D => 
                           n20, Q => n1443);
   U3591 : OAI222 port map( A => X_barycentre_top_5_port, B => n849, C => n1444
                           , D => n1443, Q => n1445);
   U3592 : OAI222 port map( A => n1446, B => n1445, C => position1_N2378, D => 
                           n25, Q => n1447);
   U3593 : OAI222 port map( A => X_barycentre_top_7_port, B => n847, C => n1448
                           , D => n1447, Q => n1449);
   U3594 : OAI222 port map( A => n1450, B => n1449, C => position1_N2380, D => 
                           n29, Q => position1_N2381);
   U3595 : OAI212 port map( A => n1452, B => n631, C => position1_n1231, Q => 
                           n1451);
   U3596 : OAI222 port map( A => position1_n1224, B => n472, C => n897, D => 
                           n896, Q => n1468);
   U3597 : OAI222 port map( A => n1468, B => n1467, C => n259, D => n895, Q => 
                           n1469);
   U3598 : OAI212 port map( A => n595, B => position1_n1264, C => n1557, Q => 
                           n1559);
   U3599 : OAI222 port map( A => n1566, B => n1565, C => n517, D => 
                           position1_n1304, Q => n1567);
   U3600 : OAI222 port map( A => n990, B => n630, C => n1568, D => n1567, Q => 
                           n1569);
   U3601 : OAI222 port map( A => n1570, B => n1569, C => n626, D => 
                           position1_n1302, Q => n1571);
   U3602 : OAI222 port map( A => n988, B => n38, C => n1572, D => n1571, Q => 
                           n1573);
   U3603 : OAI222 port map( A => n1574, B => n1573, C => n469, D => 
                           position1_n1300, Q => n1575);
   U3604 : OAI222 port map( A => n986, B => n48, C => n1576, D => n1575, Q => 
                           n1577);
   U3605 : OAI222 port map( A => n1578, B => n1577, C => n470, D => 
                           position1_n1298, Q => n1579);
   U3606 : OAI222 port map( A => n984, B => n254, C => n1580, D => n1579, Q => 
                           n1581);
   U3607 : OAI222 port map( A => n1582, B => n1581, C => n472, D => 
                           position1_n1296, Q => n1583);
   U3608 : OAI222 port map( A => n982, B => n286, C => n1584, D => n1583, Q => 
                           n1585);
   U3609 : OAI222 port map( A => n1586, B => n1585, C => n474, D => 
                           position1_n1294, Q => n1587);
   U3610 : OAI222 port map( A => n980, B => n39, C => n1588, D => n1587, Q => 
                           n1589);
   U3611 : OAI222 port map( A => n1590, B => n1589, C => n475, D => 
                           position1_n1292, Q => n1591);
   U3612 : OAI222 port map( A => n978, B => n40, C => n1592, D => n1591, Q => 
                           n1593);
   U3613 : OAI222 port map( A => n1594, B => n1593, C => n476, D => 
                           position1_n1290, Q => n1595);
   U3614 : OAI222 port map( A => n1606, B => n1021, C => n517, D => 
                           position1_n1328, Q => n1607);
   U3615 : OAI222 port map( A => n1020, B => n630, C => n1019, D => n1607, Q =>
                           n1608);
   U3616 : OAI222 port map( A => n1017, B => n1608, C => n628, D => 
                           position1_n1326, Q => n1609);
   U3617 : OAI222 port map( A => n1016, B => n38, C => n1015, D => n1609, Q => 
                           n1610);
   U3618 : OAI222 port map( A => n1013, B => n1610, C => position1_N2457, D => 
                           position1_n1324, Q => n1611);
   U3619 : OAI222 port map( A => n1011, B => n252, C => n1612, D => n1611, Q =>
                           n1613);
   U3620 : OAI212 port map( A => n633, B => n1046, C => n1641, Q => n1642);
   U3621 : OAI212 port map( A => position1_N2073, B => n630, C => n1642, Q => 
                           n1643);
   U3622 : OAI222 port map( A => n1644, B => n1643, C => n628, D => n1045, Q =>
                           n1645);
   U3623 : OAI222 port map( A => position1_N2075, B => n38, C => n1646, D => 
                           n1645, Q => n1647);
   U3624 : OAI222 port map( A => n1648, B => n1647, C => n469, D => n1043, Q =>
                           n1649);
   U3625 : OAI222 port map( A => position1_N2077, B => n48, C => n1650, D => 
                           n1649, Q => n1651);
   U3626 : OAI222 port map( A => n1652, B => n1651, C => n471, D => n1041, Q =>
                           n1653);
   U3627 : OAI222 port map( A => position1_N2079, B => n282, C => n1654, D => 
                           n1653, Q => n1655);
   U3628 : OAI222 port map( A => n1656, B => n1655, C => position1_N2453, D => 
                           n1039, Q => n1657);
   U3629 : OAI222 port map( A => position1_N2081, B => n286, C => n1658, D => 
                           n1657, Q => n1659);
   U3630 : OAI222 port map( A => n1660, B => n1659, C => n474, D => n1037, Q =>
                           n1661);
   U3631 : OAI222 port map( A => position1_N2083, B => n39, C => n1662, D => 
                           n1661, Q => n1663);
   U3632 : OAI222 port map( A => n1664, B => n1663, C => position1_N2449, D => 
                           n1035, Q => n1665);
   U3633 : OAI222 port map( A => position1_N2085, B => n40, C => n1666, D => 
                           n1665, Q => n1667);
   U3634 : OAI222 port map( A => n1668, B => n1667, C => position1_N2447, D => 
                           n1033, Q => n1669);
   U3635 : OAI222 port map( A => position1_N2087, B => n68, C => n1670, D => 
                           n1669, Q => n1671);
   U3636 : OAI222 port map( A => n1672, B => n1671, C => n595, D => n1030, Q =>
                           n1673);
   U3637 : OAI212 port map( A => n1673, B => n590, C => position1_N2089, Q => 
                           n1675);
   U3638 : OAI212 port map( A => n633, B => position1_n1350, C => n1680, Q => 
                           n1681);
   U3639 : OAI212 port map( A => n1081, B => n630, C => n1681, Q => n1682);
   U3640 : OAI222 port map( A => n1078, B => n1682, C => n628, D => 
                           position1_n1349, Q => n1683);
   U3641 : OAI222 port map( A => n1074, B => n276, C => n1684, D => n1683, Q =>
                           n1685);
   U3642 : IMAJ31 port map( A => n1083, B => n588, C => n1748, Q => 
                           position1_N1988);
   U3643 : OAI212 port map( A => n49, B => n517, C => n1349, Q => n1753);
   U3644 : OAI222 port map( A => n1753, B => n1752, C => n272, D => 
                           position1_y_sum_10_port, Q => n1754);
   U3645 : OAI212 port map( A => n1786, B => n633, C => position1_n1427, Q => 
                           n1785);
   U3646 : OAI222 port map( A => position1_n1420, B => position1_N2453, C => 
                           n1116, D => n1115, Q => n1802);
   U3647 : OAI222 port map( A => n1802, B => n1801, C => n259, D => n1114, Q =>
                           n1803);
   U3648 : OAI212 port map( A => n596, B => position1_n1460, C => n1891, Q => 
                           n1893);
   U3649 : OAI222 port map( A => n1900, B => n1899, C => n518, D => 
                           position1_n1500, Q => n1901);
   U3650 : OAI222 port map( A => n1209, B => n630, C => n1902, D => n1901, Q =>
                           n1903);
   U3651 : OAI222 port map( A => n1904, B => n1903, C => n628, D => 
                           position1_n1498, Q => n1905);
   U3652 : OAI222 port map( A => n1207, B => n38, C => n1906, D => n1905, Q => 
                           n1907);
   U3653 : OAI222 port map( A => n1908, B => n1907, C => position1_N2457, D => 
                           position1_n1496, Q => n1909);
   U3654 : OAI222 port map( A => n1205, B => n48, C => n1910, D => n1909, Q => 
                           n1911);
   U3655 : OAI222 port map( A => n1912, B => n1911, C => n470, D => 
                           position1_n1494, Q => n1913);
   U3656 : OAI222 port map( A => n1203, B => n254, C => n1914, D => n1913, Q =>
                           n1915);
   U3657 : OAI222 port map( A => n1916, B => n1915, C => n472, D => 
                           position1_n1492, Q => n1917);
   U3658 : OAI222 port map( A => n1201, B => n286, C => n1918, D => n1917, Q =>
                           n1919);
   U3659 : OAI222 port map( A => n1920, B => n1919, C => n474, D => 
                           position1_n1490, Q => n1921);
   U3660 : OAI222 port map( A => n1199, B => n39, C => n1922, D => n1921, Q => 
                           n1923);
   U3661 : OAI222 port map( A => n1924, B => n1923, C => n475, D => 
                           position1_n1488, Q => n1925);
   U3662 : OAI222 port map( A => n1197, B => n40, C => n1926, D => n1925, Q => 
                           n1927);
   U3663 : OAI222 port map( A => n1928, B => n1927, C => n476, D => 
                           position1_n1486, Q => n1929);
   U3664 : OAI222 port map( A => n1940, B => n1240, C => n518, D => 
                           position1_n1524, Q => n1941);
   U3665 : OAI222 port map( A => n1239, B => n630, C => n1238, D => n1941, Q =>
                           n1942);
   U3666 : OAI222 port map( A => n1236, B => n1942, C => n628, D => 
                           position1_n1522, Q => n1943);
   U3667 : OAI222 port map( A => n1235, B => n38, C => n1234, D => n1943, Q => 
                           n1944);
   U3668 : OAI222 port map( A => n1232, B => n1944, C => n469, D => 
                           position1_n1520, Q => n1945);
   U3669 : OAI222 port map( A => n1230, B => n46, C => n1946, D => n1945, Q => 
                           n1947);
   U3670 : OAI212 port map( A => n633, B => n1265, C => n1975, Q => n1976);
   U3671 : OAI212 port map( A => position1_N1656, B => n630, C => n1976, Q => 
                           n1977);
   U3672 : OAI222 port map( A => n1978, B => n1977, C => n628, D => n1264, Q =>
                           n1979);
   U3673 : OAI222 port map( A => position1_N1658, B => n38, C => n1980, D => 
                           n1979, Q => n1981);
   U3674 : OAI222 port map( A => n1982, B => n1981, C => position1_N2457, D => 
                           n1262, Q => n1983);
   U3675 : OAI222 port map( A => position1_N1660, B => n48, C => n1984, D => 
                           n1983, Q => n1985);
   U3676 : OAI222 port map( A => n1986, B => n1985, C => n471, D => n1260, Q =>
                           n1987);
   U3677 : OAI222 port map( A => position1_N1662, B => n101, C => n1988, D => 
                           n1987, Q => n1989);
   U3678 : OAI222 port map( A => n1990, B => n1989, C => position1_N2453, D => 
                           n1258, Q => n1991);
   U3679 : OAI222 port map( A => position1_N1664, B => n286, C => n1992, D => 
                           n1991, Q => n1993);
   U3680 : OAI222 port map( A => n1994, B => n1993, C => n474, D => n1256, Q =>
                           n1995);
   U3681 : OAI222 port map( A => position1_N1666, B => n39, C => n1996, D => 
                           n1995, Q => n1997);
   U3682 : OAI222 port map( A => n1998, B => n1997, C => position1_N2449, D => 
                           n1254, Q => n1999);
   U3683 : OAI222 port map( A => position1_N1668, B => n40, C => n2000, D => 
                           n1999, Q => n2001);
   U3684 : OAI222 port map( A => n2002, B => n2001, C => position1_N2447, D => 
                           n1252, Q => n2003);
   U3685 : OAI222 port map( A => position1_N1670, B => n68, C => n2004, D => 
                           n2003, Q => n2005);
   U3686 : OAI222 port map( A => n2006, B => n2005, C => n595, D => n1249, Q =>
                           n2007);
   U3687 : OAI212 port map( A => n2007, B => n591, C => position1_N1672, Q => 
                           n2009);
   U3688 : OAI212 port map( A => n633, B => position1_n1546, C => n2014, Q => 
                           n2015);
   U3689 : OAI212 port map( A => n1300, B => n630, C => n2015, Q => n2016);
   U3690 : OAI222 port map( A => n1297, B => n2016, C => n628, D => 
                           position1_n1545, Q => n2017);
   U3691 : OAI222 port map( A => n1293, B => n248, C => n2018, D => n2017, Q =>
                           n2019);
   U3692 : IMAJ31 port map( A => n1302, B => n588, C => n2082, Q => 
                           position1_N1571_port);
   U3693 : OAI212 port map( A => n50, B => n517, C => n1350, Q => n2087);
   U3694 : OAI222 port map( A => n2087, B => n2086, C => n67, D => 
                           position1_x_sum_10_port, Q => n2088);
   U3695 : OAI212 port map( A => n2121, B => n2120, C => n2119, Q => n2122);

end SYN_bar;
