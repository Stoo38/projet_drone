../../BENCH/test_bench.vhd