../../BENCH/bench_top_ppm.vhd