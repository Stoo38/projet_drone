../results/send_ppm.vhd