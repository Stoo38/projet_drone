../../BENCH/test_ppm.vhd