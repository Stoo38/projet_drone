
module top_bar ( CLK_top, reset_top, SW1_top, r_top, g_top, b_top, rout_top, 
        gout_top, bout_top, r_out_proc, g_out_proc, b_out_proc, 
        X_barycentre_top, Y_barycentre_top, HSYNC_top, VSYNC_top, cam_x, cam_y, 
        IMG_top );
  input [7:0] r_top;
  input [7:0] g_top;
  input [7:0] b_top;
  output [7:0] rout_top;
  output [7:0] gout_top;
  output [7:0] bout_top;
  output [7:0] r_out_proc;
  output [7:0] g_out_proc;
  output [7:0] b_out_proc;
  output [8:0] X_barycentre_top;
  output [8:0] Y_barycentre_top;
  output [9:0] cam_x;
  output [8:0] cam_y;
  input CLK_top, reset_top, SW1_top;
  output HSYNC_top, VSYNC_top, IMG_top;
  wire   \*Logic0* , n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, \gensync1/n107 , \gensync1/n106 , \gensync1/n105 ,
         \gensync1/n104 , \gensync1/n103 , \gensync1/n102 , \gensync1/n101 ,
         \gensync1/n100 , \gensync1/n99 , \gensync1/n98 , \gensync1/n97 ,
         \gensync1/n96 , \gensync1/n95 , \gensync1/n94 , \gensync1/n93 ,
         \gensync1/n92 , \gensync1/n91 , \gensync1/n90 , \gensync1/n89 ,
         \gensync1/n88 , \gensync1/n87 , \gensync1/N182 , \gensync1/N181 ,
         \gensync1/N180 , \gensync1/N179 , \gensync1/N178 , \gensync1/N177 ,
         \gensync1/N176 , \gensync1/N175 , \gensync1/N174 , \gensync1/N173 ,
         \gensync1/N172 , \gensync1/N171 , \gensync1/N170 , \gensync1/N169 ,
         \gensync1/N168 , \gensync1/N167 , \gensync1/N166 , \gensync1/N165 ,
         \gensync1/N145 , \gensync1/N144 , \gensync1/N143 , \gensync1/N142 ,
         \gensync1/N141 , \gensync1/N140 , \gensync1/N139 , \gensync1/N138 ,
         \gensync1/N135 , \gensync1/N132 , \gensync1/N129 , \gensync1/N85 ,
         \gensync1/N74 , \gensync1/N72 , \gensync1/N69 , \gensync1/N66 ,
         \gensync1/N65 , \gensync1/N64 , \gensync1/N63 , \gensync1/N62 ,
         \gensync1/N61 , \gensync1/N60 , \gensync1/N59 , \gensync1/N58 ,
         \gensync1/N57 , \gensync1/N56 , \gensync1/N54 , \gensync1/N53 ,
         \gensync1/N52 , \gensync1/N51 , \gensync1/N50 , \gensync1/N49 ,
         \gensync1/N48 , \gensync1/N47 , \gensync1/N43 , \gensync1/comptY[9] ,
         \gensync1/N31 , \gensync1/N30 , \gensync1/N29 , \gensync1/N28 ,
         \gensync1/N27 , \gensync1/N26 , \gensync1/N25 , \gensync1/N24 ,
         \gensync1/N23 , \gensync1/N22 , \gensync1/N20 , \gensync1/N19 ,
         \gensync1/N18 , \gensync1/N17 , \gensync1/N16 , \gensync1/N15 ,
         \gensync1/N14 , \gensync1/N13 , \gensync1/N9 , \image_process1/n119 ,
         \image_process1/n118 , \image_process1/n117 , \image_process1/n116 ,
         \image_process1/n115 , \image_process1/n114 , \image_process1/n113 ,
         \image_process1/n112 , \image_process1/n111 , \image_process1/n110 ,
         \image_process1/n109 , \image_process1/n108 , \image_process1/n107 ,
         \image_process1/n106 , \image_process1/n105 , \image_process1/n104 ,
         \image_process1/n103 , \image_process1/n102 , \image_process1/n101 ,
         \image_process1/n100 , \image_process1/n99 , \image_process1/n98 ,
         \image_process1/n97 , \image_process1/n96 , \image_process1/n95 ,
         \image_process1/n94 , \image_process1/n93 , \image_process1/n92 ,
         \image_process1/n91 , \image_process1/n90 , \image_process1/n89 ,
         \image_process1/n88 , \image_process1/n87 , \image_process1/n86 ,
         \image_process1/n85 , \image_process1/n84 , \image_process1/n83 ,
         \image_process1/n82 , \image_process1/n81 , \image_process1/n80 ,
         \image_process1/n79 , \image_process1/n78 , \image_process1/n77 ,
         \image_process1/n76 , \image_process1/n75 , \image_process1/n74 ,
         \image_process1/n73 , \image_process1/n72 , \image_process1/n71 ,
         \image_process1/n70 , \image_process1/n69 , \image_process1/n68 ,
         \image_process1/n67 , \image_process1/n66 , \image_process1/n65 ,
         \image_process1/n64 , \image_process1/n63 , \image_process1/n62 ,
         \image_process1/n61 , \image_process1/n60 , \image_process1/n59 ,
         \image_process1/n58 , \image_process1/n57 , \image_process1/n56 ,
         \image_process1/n55 , \image_process1/n27 , \image_process1/n25 ,
         \image_process1/n13 , \image_process1/N64 , \image_process1/N62 ,
         \image_process1/N59 , \image_process1/N31 , \image_process1/N29 ,
         \image_process1/N28 , \image_process1/N26 , \image_process1/N25 ,
         \image_process1/N23 , \image_process1/N22 , \image_process1/N20 ,
         \image_process1/N19 , \image_process1/N17 , \image_process1/N16 ,
         \image_process1/N14 , \image_process1/N13 , \image_process1/N11 ,
         \image_process1/N10 , \image_process1/N8 , \image_process1/state ,
         \position1/n1635 , \position1/n1634 , \position1/n1633 ,
         \position1/n1632 , \position1/n1631 , \position1/n1630 ,
         \position1/n1629 , \position1/n1628 , \position1/n1627 ,
         \position1/n1626 , \position1/n1625 , \position1/n1624 ,
         \position1/n1623 , \position1/n1622 , \position1/n1621 ,
         \position1/n1620 , \position1/n1619 , \position1/n1618 ,
         \position1/n1617 , \position1/n1616 , \position1/n1615 ,
         \position1/n1614 , \position1/n1613 , \position1/n1612 ,
         \position1/n1611 , \position1/n1610 , \position1/n1609 ,
         \position1/n1608 , \position1/n1607 , \position1/n1606 ,
         \position1/n1605 , \position1/n1604 , \position1/n1603 ,
         \position1/n1602 , \position1/n1601 , \position1/n1600 ,
         \position1/n1599 , \position1/n1598 , \position1/n1597 ,
         \position1/n1596 , \position1/n1595 , \position1/n1594 ,
         \position1/n1593 , \position1/n1592 , \position1/n1591 ,
         \position1/n1590 , \position1/n1589 , \position1/n1588 ,
         \position1/n1587 , \position1/n1586 , \position1/n1585 ,
         \position1/n1584 , \position1/n1583 , \position1/n1582 ,
         \position1/n1581 , \position1/n1580 , \position1/n1579 ,
         \position1/n1578 , \position1/n1577 , \position1/n1576 ,
         \position1/n1575 , \position1/n1574 , \position1/n1573 ,
         \position1/n1572 , \position1/n1571 , \position1/n1570 ,
         \position1/n1569 , \position1/n1568 , \position1/n1567 ,
         \position1/n1566 , \position1/n1565 , \position1/n1564 ,
         \position1/n1563 , \position1/n1562 , \position1/n1561 ,
         \position1/n1560 , \position1/n1559 , \position1/n1558 ,
         \position1/n1557 , \position1/n1556 , \position1/n1555 ,
         \position1/n1554 , \position1/n1553 , \position1/n1552 ,
         \position1/n1551 , \position1/n1550 , \position1/n1549 ,
         \position1/n1548 , \position1/n1547 , \position1/n1546 ,
         \position1/n1545 , \position1/n1544 , \position1/n1543 ,
         \position1/n1542 , \position1/n1541 , \position1/n1540 ,
         \position1/n1539 , \position1/n1538 , \position1/n1537 ,
         \position1/n1536 , \position1/n1535 , \position1/n1534 ,
         \position1/n1533 , \position1/n1532 , \position1/n1531 ,
         \position1/n1530 , \position1/n1529 , \position1/n1528 ,
         \position1/n1527 , \position1/n1526 , \position1/n1525 ,
         \position1/n1524 , \position1/n1523 , \position1/n1522 ,
         \position1/n1521 , \position1/n1520 , \position1/n1519 ,
         \position1/n1518 , \position1/n1517 , \position1/n1516 ,
         \position1/n1515 , \position1/n1514 , \position1/n1513 ,
         \position1/n1512 , \position1/n1511 , \position1/n1510 ,
         \position1/n1509 , \position1/n1508 , \position1/n1507 ,
         \position1/n1506 , \position1/n1505 , \position1/n1504 ,
         \position1/n1503 , \position1/n1502 , \position1/n1501 ,
         \position1/n1500 , \position1/n1499 , \position1/n1498 ,
         \position1/n1497 , \position1/n1496 , \position1/n1495 ,
         \position1/n1494 , \position1/n1493 , \position1/n1492 ,
         \position1/n1491 , \position1/n1490 , \position1/n1489 ,
         \position1/n1488 , \position1/n1487 , \position1/n1486 ,
         \position1/n1485 , \position1/n1484 , \position1/n1483 ,
         \position1/n1482 , \position1/n1481 , \position1/n1480 ,
         \position1/n1479 , \position1/n1478 , \position1/n1477 ,
         \position1/n1476 , \position1/n1475 , \position1/n1474 ,
         \position1/n1473 , \position1/n1472 , \position1/n1471 ,
         \position1/n1470 , \position1/n1469 , \position1/n1468 ,
         \position1/n1467 , \position1/n1466 , \position1/n1465 ,
         \position1/n1464 , \position1/n1463 , \position1/n1462 ,
         \position1/n1461 , \position1/n1460 , \position1/n1459 ,
         \position1/n1458 , \position1/n1457 , \position1/n1456 ,
         \position1/n1455 , \position1/n1454 , \position1/n1453 ,
         \position1/n1452 , \position1/n1451 , \position1/n1450 ,
         \position1/n1449 , \position1/n1448 , \position1/n1447 ,
         \position1/n1446 , \position1/n1445 , \position1/n1444 ,
         \position1/n1443 , \position1/n1442 , \position1/n1441 ,
         \position1/n1440 , \position1/n1439 , \position1/n1438 ,
         \position1/n1437 , \position1/n1436 , \position1/n1435 ,
         \position1/n1434 , \position1/n1433 , \position1/n1432 ,
         \position1/n1431 , \position1/n1430 , \position1/n1429 ,
         \position1/n1428 , \position1/n1427 , \position1/n1426 ,
         \position1/n1425 , \position1/n1424 , \position1/n1423 ,
         \position1/n1422 , \position1/n1421 , \position1/n1420 ,
         \position1/n1419 , \position1/n1418 , \position1/n1417 ,
         \position1/n1416 , \position1/n1415 , \position1/n1414 ,
         \position1/n1413 , \position1/n1412 , \position1/n1411 ,
         \position1/n1410 , \position1/n1409 , \position1/n1408 ,
         \position1/n1407 , \position1/n1406 , \position1/n1405 ,
         \position1/n1404 , \position1/n1403 , \position1/n1402 ,
         \position1/n1401 , \position1/n1400 , \position1/n1399 ,
         \position1/n1398 , \position1/n1397 , \position1/n1396 ,
         \position1/n1395 , \position1/n1394 , \position1/n1393 ,
         \position1/n1392 , \position1/n1391 , \position1/n1390 ,
         \position1/n1389 , \position1/n1388 , \position1/n1387 ,
         \position1/n1386 , \position1/n1385 , \position1/n1384 ,
         \position1/n1383 , \position1/n1382 , \position1/n1381 ,
         \position1/n1380 , \position1/n1379 , \position1/n1378 ,
         \position1/n1377 , \position1/n1376 , \position1/n1375 ,
         \position1/n1374 , \position1/n1373 , \position1/n1372 ,
         \position1/n1371 , \position1/n1370 , \position1/n1369 ,
         \position1/n1368 , \position1/n1367 , \position1/n1366 ,
         \position1/n1365 , \position1/n1364 , \position1/n1363 ,
         \position1/n1362 , \position1/n1361 , \position1/n1360 ,
         \position1/n1359 , \position1/n1358 , \position1/n1357 ,
         \position1/n1356 , \position1/n1355 , \position1/n1354 ,
         \position1/n1353 , \position1/n1352 , \position1/n1351 ,
         \position1/n1350 , \position1/n1349 , \position1/n1348 ,
         \position1/n1347 , \position1/n1346 , \position1/n1345 ,
         \position1/n1344 , \position1/n1343 , \position1/n1342 ,
         \position1/n1341 , \position1/n1340 , \position1/n1339 ,
         \position1/n1338 , \position1/n1337 , \position1/n1336 ,
         \position1/n1335 , \position1/n1334 , \position1/n1333 ,
         \position1/n1332 , \position1/n1331 , \position1/n1330 ,
         \position1/n1329 , \position1/n1328 , \position1/n1327 ,
         \position1/n1326 , \position1/n1325 , \position1/n1324 ,
         \position1/n1323 , \position1/n1322 , \position1/n1321 ,
         \position1/n1320 , \position1/n1319 , \position1/n1318 ,
         \position1/n1317 , \position1/n1316 , \position1/n1315 ,
         \position1/n1314 , \position1/n1313 , \position1/n1312 ,
         \position1/n1311 , \position1/n1310 , \position1/n1309 ,
         \position1/n1308 , \position1/n1307 , \position1/n1306 ,
         \position1/n1305 , \position1/n1304 , \position1/n1303 ,
         \position1/n1302 , \position1/n1301 , \position1/n1300 ,
         \position1/n1299 , \position1/n1298 , \position1/n1297 ,
         \position1/n1296 , \position1/n1295 , \position1/n1294 ,
         \position1/n1293 , \position1/n1292 , \position1/n1291 ,
         \position1/n1290 , \position1/n1289 , \position1/n1288 ,
         \position1/n1287 , \position1/n1286 , \position1/n1285 ,
         \position1/n1284 , \position1/n1283 , \position1/n1282 ,
         \position1/n1281 , \position1/n1280 , \position1/n1279 ,
         \position1/n1278 , \position1/n1277 , \position1/n1276 ,
         \position1/n1275 , \position1/n1274 , \position1/n1273 ,
         \position1/n1272 , \position1/n1271 , \position1/n1270 ,
         \position1/n1269 , \position1/n1268 , \position1/n1267 ,
         \position1/n1266 , \position1/n1265 , \position1/n1264 ,
         \position1/n1263 , \position1/n1262 , \position1/n1261 ,
         \position1/n1260 , \position1/n1259 , \position1/n1258 ,
         \position1/n1257 , \position1/n1256 , \position1/n1255 ,
         \position1/n1254 , \position1/n1253 , \position1/n1252 ,
         \position1/n1251 , \position1/n1250 , \position1/n1249 ,
         \position1/n1248 , \position1/n1247 , \position1/n1246 ,
         \position1/n1245 , \position1/n1244 , \position1/n1243 ,
         \position1/n1242 , \position1/n1241 , \position1/n1240 ,
         \position1/n1239 , \position1/n1238 , \position1/n1237 ,
         \position1/n1236 , \position1/n1235 , \position1/n1234 ,
         \position1/n1233 , \position1/n1232 , \position1/n1231 ,
         \position1/n1230 , \position1/n1229 , \position1/n1228 ,
         \position1/n1227 , \position1/n1226 , \position1/n1225 ,
         \position1/n1224 , \position1/n1223 , \position1/n1222 ,
         \position1/n1221 , \position1/n1220 , \position1/n1219 ,
         \position1/n1218 , \position1/n1217 , \position1/n1216 ,
         \position1/n1215 , \position1/n1214 , \position1/n1213 ,
         \position1/n1212 , \position1/n1211 , \position1/n1210 ,
         \position1/n1209 , \position1/n1208 , \position1/n1207 ,
         \position1/n1206 , \position1/n1205 , \position1/n1204 ,
         \position1/n1203 , \position1/n1202 , \position1/n1201 ,
         \position1/n1200 , \position1/n1199 , \position1/n1198 ,
         \position1/n1197 , \position1/n1196 , \position1/n1195 ,
         \position1/n1194 , \position1/n1193 , \position1/n1192 ,
         \position1/n1191 , \position1/n1190 , \position1/n1189 ,
         \position1/n1188 , \position1/n1187 , \position1/n1186 ,
         \position1/n1185 , \position1/n1184 , \position1/n1183 ,
         \position1/n1182 , \position1/n1181 , \position1/n1180 ,
         \position1/n1179 , \position1/n1178 , \position1/n1177 ,
         \position1/n1176 , \position1/n1175 , \position1/n1174 ,
         \position1/n1173 , \position1/n1172 , \position1/n1171 ,
         \position1/n1170 , \position1/n1169 , \position1/n1168 ,
         \position1/n1167 , \position1/n1166 , \position1/n1165 ,
         \position1/n1164 , \position1/n1163 , \position1/n1162 ,
         \position1/n1161 , \position1/n1160 , \position1/n1159 ,
         \position1/n1158 , \position1/n1157 , \position1/n1156 ,
         \position1/n1154 , \position1/n1153 , \position1/n1152 ,
         \position1/n1151 , \position1/n1150 , \position1/n1149 ,
         \position1/n1148 , \position1/n1147 , \position1/n1146 ,
         \position1/n1145 , \position1/n1144 , \position1/n1143 ,
         \position1/n1142 , \position1/n1141 , \position1/n1140 ,
         \position1/n1139 , \position1/n1138 , \position1/n1137 ,
         \position1/n1136 , \position1/n1135 , \position1/n1134 ,
         \position1/n1133 , \position1/n1132 , \position1/n1131 ,
         \position1/n1130 , \position1/n1129 , \position1/n1128 ,
         \position1/n1127 , \position1/n1126 , \position1/n1125 ,
         \position1/n1124 , \position1/n1123 , \position1/n1122 ,
         \position1/n1121 , \position1/n1120 , \position1/n1119 ,
         \position1/n1118 , \position1/n1117 , \position1/n1116 ,
         \position1/n1115 , \position1/n1114 , \position1/n1113 ,
         \position1/n1112 , \position1/n1111 , \position1/n1110 ,
         \position1/n1109 , \position1/n1108 , \position1/n1107 ,
         \position1/n1106 , \position1/n1105 , \position1/n1104 ,
         \position1/n1103 , \position1/n1102 , \position1/n1101 ,
         \position1/n1100 , \position1/n1099 , \position1/n1098 ,
         \position1/n1097 , \position1/n1096 , \position1/n1095 ,
         \position1/n1094 , \position1/n1093 , \position1/n1092 ,
         \position1/n1091 , \position1/n1090 , \position1/n1089 ,
         \position1/n1088 , \position1/n1087 , \position1/n1086 ,
         \position1/n1085 , \position1/n1084 , \position1/n1083 ,
         \position1/n1082 , \position1/n1081 , \position1/n1080 ,
         \position1/n1079 , \position1/n1078 , \position1/n1077 ,
         \position1/n1076 , \position1/n1075 , \position1/n1074 ,
         \position1/n1073 , \position1/n1072 , \position1/n1071 ,
         \position1/n1070 , \position1/n1069 , \position1/n1068 ,
         \position1/n1067 , \position1/n1066 , \position1/n1065 ,
         \position1/n1064 , \position1/n1063 , \position1/n1062 ,
         \position1/n1061 , \position1/n1060 , \position1/n1059 ,
         \position1/n1058 , \position1/n1057 , \position1/n1056 ,
         \position1/n1055 , \position1/n1054 , \position1/n1053 ,
         \position1/n1052 , \position1/n1051 , \position1/n1050 ,
         \position1/n1049 , \position1/n1048 , \position1/n1047 ,
         \position1/n1046 , \position1/n1045 , \position1/n1044 ,
         \position1/n1043 , \position1/n1042 , \position1/n1041 ,
         \position1/n1040 , \position1/n1039 , \position1/n1038 ,
         \position1/n1037 , \position1/n1036 , \position1/n1035 ,
         \position1/n1034 , \position1/n1033 , \position1/n1032 ,
         \position1/n1031 , \position1/n1030 , \position1/n1029 ,
         \position1/n1028 , \position1/n1027 , \position1/n1026 ,
         \position1/n1025 , \position1/n1024 , \position1/n1023 ,
         \position1/n1022 , \position1/n1021 , \position1/n1020 ,
         \position1/n1019 , \position1/n1018 , \position1/n1017 ,
         \position1/n1016 , \position1/n1015 , \position1/n1014 ,
         \position1/n1013 , \position1/n1012 , \position1/n1011 ,
         \position1/n1010 , \position1/n1009 , \position1/n1008 ,
         \position1/n1007 , \position1/n1006 , \position1/n1005 ,
         \position1/n1004 , \position1/n1003 , \position1/n1002 ,
         \position1/n1001 , \position1/n1000 , \position1/n999 ,
         \position1/n998 , \position1/n997 , \position1/n996 ,
         \position1/n995 , \position1/n994 , \position1/n993 ,
         \position1/n992 , \position1/n991 , \position1/n990 ,
         \position1/n989 , \position1/n988 , \position1/n987 ,
         \position1/n986 , \position1/n985 , \position1/n984 ,
         \position1/n983 , \position1/n982 , \position1/n981 ,
         \position1/n980 , \position1/n979 , \position1/n978 ,
         \position1/n977 , \position1/n976 , \position1/n975 ,
         \position1/n974 , \position1/n973 , \position1/n972 ,
         \position1/n971 , \position1/n970 , \position1/n969 ,
         \position1/n968 , \position1/n967 , \position1/n966 ,
         \position1/n965 , \position1/n964 , \position1/n963 ,
         \position1/n962 , \position1/n961 , \position1/n960 ,
         \position1/n959 , \position1/n958 , \position1/n957 ,
         \position1/n956 , \position1/n955 , \position1/n954 ,
         \position1/n953 , \position1/n952 , \position1/n951 ,
         \position1/n950 , \position1/n949 , \position1/n948 ,
         \position1/n947 , \position1/n946 , \position1/n945 ,
         \position1/n944 , \position1/n943 , \position1/n942 ,
         \position1/n941 , \position1/n940 , \position1/n939 ,
         \position1/n938 , \position1/n937 , \position1/n936 ,
         \position1/n935 , \position1/n934 , \position1/n933 ,
         \position1/n932 , \position1/n931 , \position1/n930 ,
         \position1/n929 , \position1/n928 , \position1/n927 ,
         \position1/n926 , \position1/n925 , \position1/n924 ,
         \position1/n923 , \position1/n922 , \position1/n921 ,
         \position1/n920 , \position1/n919 , \position1/n918 ,
         \position1/n917 , \position1/n916 , \position1/n915 ,
         \position1/n914 , \position1/n913 , \position1/n912 ,
         \position1/n911 , \position1/n910 , \position1/n909 ,
         \position1/n908 , \position1/n907 , \position1/n906 ,
         \position1/n905 , \position1/n904 , \position1/n903 ,
         \position1/n902 , \position1/n901 , \position1/n900 ,
         \position1/n899 , \position1/n898 , \position1/n897 ,
         \position1/n896 , \position1/n895 , \position1/n894 ,
         \position1/n893 , \position1/n892 , \position1/n891 ,
         \position1/n890 , \position1/n889 , \position1/n888 ,
         \position1/n887 , \position1/n886 , \position1/n885 ,
         \position1/n884 , \position1/n883 , \position1/n882 ,
         \position1/n881 , \position1/n880 , \position1/n879 ,
         \position1/n878 , \position1/n877 , \position1/n876 ,
         \position1/n875 , \position1/n874 , \position1/n873 ,
         \position1/n872 , \position1/n871 , \position1/n870 ,
         \position1/n869 , \position1/n868 , \position1/n867 ,
         \position1/n866 , \position1/n865 , \position1/n864 ,
         \position1/n863 , \position1/n862 , \position1/n861 ,
         \position1/n860 , \position1/n859 , \position1/n858 ,
         \position1/n857 , \position1/n856 , \position1/n855 ,
         \position1/n854 , \position1/n853 , \position1/n852 ,
         \position1/n851 , \position1/n850 , \position1/n849 ,
         \position1/n848 , \position1/n847 , \position1/n846 ,
         \position1/n845 , \position1/n844 , \position1/n843 ,
         \position1/n842 , \position1/n841 , \position1/n840 ,
         \position1/n839 , \position1/n838 , \position1/n837 ,
         \position1/n836 , \position1/n835 , \position1/n834 ,
         \position1/n833 , \position1/n802 , \position1/n370 ,
         \position1/n369 , \position1/n368 , \position1/n367 ,
         \position1/n366 , \position1/n365 , \position1/n364 ,
         \position1/n363 , \position1/n362 , \position1/n360 ,
         \position1/n358 , \position1/n357 , \position1/n356 ,
         \position1/n353 , \position1/n352 , \position1/n351 ,
         \position1/n350 , \position1/n349 , \position1/n348 ,
         \position1/n347 , \position1/n346 , \position1/n344 ,
         \position1/n283 , \position1/dp_cluster_7/N314 ,
         \position1/dp_cluster_6/N389 , \position1/N2460 , \position1/N2459 ,
         \position1/N2458 , \position1/N2457 , \position1/N2456 ,
         \position1/N2455 , \position1/N2454 , \position1/N2453 ,
         \position1/N2452 , \position1/N2451 , \position1/N2450 ,
         \position1/N2449 , \position1/N2448 , \position1/N2447 ,
         \position1/N2446 , \position1/N2445 , \position1/N2413 ,
         \position1/N2412 , \position1/N2411 , \position1/N2410 ,
         \position1/N2409 , \position1/N2408 , \position1/N2407 ,
         \position1/N2406 , \position1/N2405 , \position1/N2402 ,
         \position1/N2401 , \position1/N2400 , \position1/N2399 ,
         \position1/N2398 , \position1/N2397 , \position1/N2396 ,
         \position1/N2395 , \position1/N2394 , \position1/N2391 ,
         \position1/N2390 , \position1/N2389 , \position1/N2388 ,
         \position1/N2387 , \position1/N2386 , \position1/N2385 ,
         \position1/N2384 , \position1/N2383 , \position1/N2381 ,
         \position1/N2380 , \position1/N2379 , \position1/N2378 ,
         \position1/N2377 , \position1/N2376 , \position1/N2375 ,
         \position1/N2374 , \position1/N2373 , \position1/N2371 ,
         \position1/N2370 , \position1/N2369 , \position1/N2368 ,
         \position1/N2367 , \position1/N2366 , \position1/N2365 ,
         \position1/N2364 , \position1/N2363 , \position1/N2362 ,
         \position1/N2361 , \position1/N2360 , \position1/N2359 ,
         \position1/N2358 , \position1/N2357 , \position1/N2356 ,
         \position1/N2355 , \position1/N2354 , \position1/N2353 ,
         \position1/N2352 , \position1/N2326 , \position1/N2325 ,
         \position1/N2324 , \position1/N2323 , \position1/N2322 ,
         \position1/N2321 , \position1/N2320 , \position1/N2319 ,
         \position1/N2318 , \position1/N2317 , \position1/N2316 ,
         \position1/N2315 , \position1/N2314 , \position1/N2313 ,
         \position1/N2312 , \position1/N2311 , \position1/N2310 ,
         \position1/N2309 , \position1/N2308 , \position1/N2307 ,
         \position1/N2306 , \position1/N2305 , \position1/N2304 ,
         \position1/N2303 , \position1/N2300 , \position1/N2274 ,
         \position1/N2273 , \position1/N2272 , \position1/N2271 ,
         \position1/N2270 , \position1/N2269 , \position1/N2268 ,
         \position1/N2267 , \position1/N2266 , \position1/N2265 ,
         \position1/N2264 , \position1/N2263 , \position1/N2262 ,
         \position1/N2261 , \position1/N2260 , \position1/N2259 ,
         \position1/N2258 , \position1/N2257 , \position1/N2256 ,
         \position1/N2255 , \position1/N2254 , \position1/N2253 ,
         \position1/N2252 , \position1/N2248 , \position1/N2222 ,
         \position1/N2221 , \position1/N2220 , \position1/N2219 ,
         \position1/N2218 , \position1/N2217 , \position1/N2216 ,
         \position1/N2215 , \position1/N2214 , \position1/N2213 ,
         \position1/N2212 , \position1/N2211 , \position1/N2210 ,
         \position1/N2209 , \position1/N2208 , \position1/N2207 ,
         \position1/N2206 , \position1/N2205 , \position1/N2204 ,
         \position1/N2203 , \position1/N2202 , \position1/N2201 ,
         \position1/N2196 , \position1/N2170 , \position1/N2169 ,
         \position1/N2168 , \position1/N2167 , \position1/N2166 ,
         \position1/N2165 , \position1/N2164 , \position1/N2163 ,
         \position1/N2162 , \position1/N2161 , \position1/N2160 ,
         \position1/N2159 , \position1/N2158 , \position1/N2157 ,
         \position1/N2156 , \position1/N2155 , \position1/N2154 ,
         \position1/N2153 , \position1/N2152 , \position1/N2151 ,
         \position1/N2150 , \position1/N2144 , \position1/N2118 ,
         \position1/N2117 , \position1/N2116 , \position1/N2115 ,
         \position1/N2114 , \position1/N2113 , \position1/N2112 ,
         \position1/N2111 , \position1/N2110 , \position1/N2109 ,
         \position1/N2108 , \position1/N2107 , \position1/N2106 ,
         \position1/N2105 , \position1/N2104 , \position1/N2103 ,
         \position1/N2102 , \position1/N2101 , \position1/N2100 ,
         \position1/N2099 , \position1/N2094 , \position1/N2092 ,
         \position1/N2091 , \position1/N2090 , \position1/N2089 ,
         \position1/N2088 , \position1/N2087 , \position1/N2086 ,
         \position1/N2085 , \position1/N2084 , \position1/N2083 ,
         \position1/N2082 , \position1/N2081 , \position1/N2080 ,
         \position1/N2079 , \position1/N2078 , \position1/N2077 ,
         \position1/N2076 , \position1/N2075 , \position1/N2074 ,
         \position1/N2073 , \position1/N2072 , \position1/N2071 ,
         \position1/N2070 , \position1/N2069 , \position1/N2068 ,
         \position1/N2065 , \position1/N2064 , \position1/N2063 ,
         \position1/N2062 , \position1/N2061 , \position1/N2060 ,
         \position1/N2059 , \position1/N2058 , \position1/N2057 ,
         \position1/N2056 , \position1/N2055 , \position1/N2054 ,
         \position1/N2053 , \position1/N2052 , \position1/N2051 ,
         \position1/N2050 , \position1/N2049 , \position1/N2040 ,
         \position1/N2014 , \position1/N2013 , \position1/N2012 ,
         \position1/N2011 , \position1/N2010 , \position1/N2009 ,
         \position1/N2008 , \position1/N2007 , \position1/N2006 ,
         \position1/N2005 , \position1/N2004 , \position1/N2003 ,
         \position1/N2002 , \position1/N2001 , \position1/N2000 ,
         \position1/N1999 , \position1/N1998 , \position1/N1997 ,
         \position1/N1990 , \position1/N1988 , \position1/N1987 ,
         \position1/N1986 , \position1/N1985 , \position1/N1984 ,
         \position1/N1983 , \position1/N1982 , \position1/N1981 ,
         \position1/N1980 , \position1/N1979 , \position1/N1978 ,
         \position1/N1977 , \position1/N1976 , \position1/N1975 ,
         \position1/N1974 , \position1/N1973 , \position1/N1972 ,
         \position1/N1971 , \position1/N1970 , \position1/N1969 ,
         \position1/N1968 , \position1/N1967 , \position1/N1966 ,
         \position1/N1965 , \position1/N1964 , \position1/N1962 ,
         \position1/N1961 , \position1/N1960 , \position1/N1959 ,
         \position1/N1958 , \position1/N1957 , \position1/N1956 ,
         \position1/N1955 , \position1/N1954 , \position1/N1953 ,
         \position1/N1952 , \position1/N1951 , \position1/N1950 ,
         \position1/N1949 , \position1/N1948 , \position1/N1947 ,
         \position1/N1946 , \position1/N1938 , \position1/N1936 ,
         \position1/N1935 , \position1/N1909 , \position1/N1908 ,
         \position1/N1907 , \position1/N1906 , \position1/N1905 ,
         \position1/N1904 , \position1/N1903 , \position1/N1902 ,
         \position1/N1901 , \position1/N1900 , \position1/N1899 ,
         \position1/N1898 , \position1/N1897 , \position1/N1896 ,
         \position1/N1895 , \position1/N1894 , \position1/N1893 ,
         \position1/N1892 , \position1/N1891 , \position1/N1890 ,
         \position1/N1889 , \position1/N1888 , \position1/N1887 ,
         \position1/N1886 , \position1/N1883 , \position1/N1857 ,
         \position1/N1856 , \position1/N1855 , \position1/N1854 ,
         \position1/N1853 , \position1/N1852 , \position1/N1851 ,
         \position1/N1850 , \position1/N1849 , \position1/N1848 ,
         \position1/N1847 , \position1/N1846 , \position1/N1845 ,
         \position1/N1844 , \position1/N1843 , \position1/N1842 ,
         \position1/N1841 , \position1/N1840 , \position1/N1839 ,
         \position1/N1838 , \position1/N1837 , \position1/N1836 ,
         \position1/N1835 , \position1/N1831 , \position1/N1805 ,
         \position1/N1804 , \position1/N1803 , \position1/N1802 ,
         \position1/N1801 , \position1/N1800 , \position1/N1799 ,
         \position1/N1798 , \position1/N1797 , \position1/N1796 ,
         \position1/N1795 , \position1/N1794 , \position1/N1793 ,
         \position1/N1792 , \position1/N1791 , \position1/N1790 ,
         \position1/N1789 , \position1/N1788 , \position1/N1787 ,
         \position1/N1786 , \position1/N1785 , \position1/N1784 ,
         \position1/N1779 , \position1/N1753 , \position1/N1752 ,
         \position1/N1751 , \position1/N1750 , \position1/N1749 ,
         \position1/N1748 , \position1/N1747 , \position1/N1746 ,
         \position1/N1745 , \position1/N1744 , \position1/N1743 ,
         \position1/N1742 , \position1/N1741 , \position1/N1740 ,
         \position1/N1739 , \position1/N1738 , \position1/N1737 ,
         \position1/N1736 , \position1/N1735 , \position1/N1734 ,
         \position1/N1733 , \position1/N1727 , \position1/N1701 ,
         \position1/N1700 , \position1/N1699 , \position1/N1698 ,
         \position1/N1697 , \position1/N1696 , \position1/N1695 ,
         \position1/N1694 , \position1/N1693 , \position1/N1692 ,
         \position1/N1691 , \position1/N1690 , \position1/N1689 ,
         \position1/N1688 , \position1/N1687 , \position1/N1686 ,
         \position1/N1685 , \position1/N1684 , \position1/N1683 ,
         \position1/N1682 , \position1/N1677 , \position1/N1675 ,
         \position1/N1674 , \position1/N1673 , \position1/N1672 ,
         \position1/N1671 , \position1/N1670 , \position1/N1669 ,
         \position1/N1668 , \position1/N1667 , \position1/N1666 ,
         \position1/N1665 , \position1/N1664 , \position1/N1663 ,
         \position1/N1662 , \position1/N1661 , \position1/N1660 ,
         \position1/N1659 , \position1/N1658 , \position1/N1657 ,
         \position1/N1656 , \position1/N1655 , \position1/N1654 ,
         \position1/N1653 , \position1/N1652 , \position1/N1651 ,
         \position1/N1648 , \position1/N1647 , \position1/N1646 ,
         \position1/N1645 , \position1/N1644 , \position1/N1643 ,
         \position1/N1642 , \position1/N1641 , \position1/N1640 ,
         \position1/N1639 , \position1/N1638 , \position1/N1637 ,
         \position1/N1636 , \position1/N1635 , \position1/N1634 ,
         \position1/N1633 , \position1/N1632 , \position1/N1623 ,
         \position1/N1597 , \position1/N1596 , \position1/N1595 ,
         \position1/N1594 , \position1/N1593 , \position1/N1592 ,
         \position1/N1591 , \position1/N1590 , \position1/N1589 ,
         \position1/N1588 , \position1/N1587 , \position1/N1586 ,
         \position1/N1585 , \position1/N1584 , \position1/N1583 ,
         \position1/N1582 , \position1/N1581 , \position1/N1580 ,
         \position1/N1573 , \position1/N1571 , \position1/N1570 ,
         \position1/N1569 , \position1/N1568 , \position1/N1567 ,
         \position1/N1566 , \position1/N1565 , \position1/N1564 ,
         \position1/N1563 , \position1/N1562 , \position1/N1561 ,
         \position1/N1560 , \position1/N1559 , \position1/N1558 ,
         \position1/N1557 , \position1/N1556 , \position1/N1555 ,
         \position1/N1554 , \position1/N1553 , \position1/N1552 ,
         \position1/N1551 , \position1/N1550 , \position1/N1549 ,
         \position1/N1548 , \position1/N1547 , \position1/N1545 ,
         \position1/N1544 , \position1/N1543 , \position1/N1542 ,
         \position1/N1541 , \position1/N1540 , \position1/N1539 ,
         \position1/N1538 , \position1/N1537 , \position1/N1536 ,
         \position1/N1535 , \position1/N1534 , \position1/N1533 ,
         \position1/N1532 , \position1/N1531 , \position1/N1530 ,
         \position1/N1529 , \position1/N1521 , \position1/N1519 ,
         \position1/N1226 , \position1/N1225 , \position1/N1224 ,
         \position1/N1223 , \position1/N1222 , \position1/N1221 ,
         \position1/N1220 , \position1/N1219 , \position1/N1218 ,
         \position1/N1217 , \position1/N1216 , \position1/N1215 ,
         \position1/N1214 , \position1/N1213 , \position1/N1212 ,
         \position1/N1211 , \position1/N1210 , \position1/N1209 ,
         \position1/N1208 , \position1/N1207 , \position1/N1206 ,
         \position1/N1205 , \position1/N1204 , \position1/N1203 ,
         \position1/N1202 , \position1/N1201 , \position1/N1200 ,
         \position1/N1199 , \position1/N1198 , \position1/N1197 ,
         \position1/N1196 , \position1/N1195 , \position1/N1194 ,
         \position1/N1193 , \position1/N1192 , \position1/N1191 ,
         \position1/N1190 , \position1/N1189 , \position1/N1188 ,
         \position1/N1187 , \position1/N1186 , \position1/N1185 ,
         \position1/N1184 , \position1/N1183 , \position1/N1182 ,
         \position1/N1181 , \position1/N1180 , \position1/N1179 ,
         \position1/N1178 , \position1/N1177 , \position1/N1003 ,
         \position1/N1002 , \position1/N1001 , \position1/N1000 ,
         \position1/N999 , \position1/N998 , \position1/N997 ,
         \position1/N996 , \position1/N995 , \position1/N994 ,
         \position1/N993 , \position1/N992 , \position1/N991 ,
         \position1/N990 , \position1/N989 , \position1/N988 ,
         \position1/N987 , \position1/N986 , \position1/N985 ,
         \position1/N984 , \position1/N983 , \position1/N982 ,
         \position1/N981 , \position1/N980 , \position1/N928 ,
         \position1/N927 , \position1/N926 , \position1/N925 ,
         \position1/N924 , \position1/N923 , \position1/N922 ,
         \position1/N921 , \position1/N920 , \position1/N919 ,
         \position1/N918 , \position1/N917 , \position1/N916 ,
         \position1/N915 , \position1/N914 , \position1/N913 ,
         \position1/N912 , \position1/N911 , \position1/N910 ,
         \position1/N909 , \position1/N908 , \position1/N907 ,
         \position1/N906 , \position1/N905 , \position1/N656 ,
         \position1/N655 , \position1/N654 , \position1/N653 ,
         \position1/N652 , \position1/N651 , \position1/N650 ,
         \position1/N649 , \position1/N648 , \position1/N647 ,
         \position1/N646 , \position1/N645 , \position1/N644 ,
         \position1/N643 , \position1/N642 , \position1/N641 ,
         \position1/N640 , \position1/N639 , \position1/N638 ,
         \position1/N637 , \position1/N636 , \position1/N635 ,
         \position1/N634 , \position1/N633 , \position1/N632 ,
         \position1/N631 , \position1/N630 , \position1/N629 ,
         \position1/N628 , \position1/N627 , \position1/N626 ,
         \position1/N625 , \position1/N624 , \position1/N623 ,
         \position1/N622 , \position1/N621 , \position1/N620 ,
         \position1/N619 , \position1/N618 , \position1/N617 ,
         \position1/N616 , \position1/N615 , \position1/N614 ,
         \position1/N613 , \position1/N612 , \position1/N611 ,
         \position1/N610 , \position1/N609 , \position1/N608 ,
         \position1/N607 , \position1/N606 , \position1/N605 ,
         \position1/N604 , \position1/N603 , \position1/N602 ,
         \position1/N601 , \position1/N600 , \position1/N599 ,
         \position1/N598 , \position1/N597 , \position1/N596 ,
         \position1/N595 , \position1/N594 , \position1/N593 ,
         \position1/N592 , \position1/N591 , \position1/N590 ,
         \position1/N577 , \position1/N576 , \position1/N575 ,
         \position1/N574 , \position1/N573 , \position1/N572 ,
         \position1/N571 , \position1/N570 , \position1/N569 ,
         \position1/N568 , \position1/N567 , \position1/N566 ,
         \position1/N565 , \position1/N564 , \position1/N563 ,
         \position1/N562 , \position1/N560 , \position1/N559 ,
         \position1/N558 , \position1/N557 , \position1/N556 ,
         \position1/N555 , \position1/N554 , \position1/N553 ,
         \position1/N552 , \position1/N551 , \position1/N550 ,
         \position1/N549 , \position1/N548 , \position1/N547 ,
         \position1/N546 , \position1/N545 , \position1/N544 ,
         \position1/N543 , \position1/N542 , \position1/N541 ,
         \position1/N540 , \position1/N539 , \position1/N538 ,
         \position1/N537 , \position1/N536 , \position1/N535 ,
         \position1/N509 , \position1/N508 , \position1/N507 ,
         \position1/N506 , \position1/N505 , \position1/N504 ,
         \position1/N503 , \position1/N502 , \position1/N501 ,
         \position1/N500 , \position1/N499 , \position1/N498 ,
         \position1/N497 , \position1/N496 , \position1/N495 ,
         \position1/N494 , \position1/N493 , \position1/N492 ,
         \position1/N491 , \position1/N490 , \position1/N489 ,
         \position1/N488 , \position1/N487 , \position1/N486 ,
         \position1/N485 , \position1/N447 , \position1/N446 ,
         \position1/N445 , \position1/N444 , \position1/N443 ,
         \position1/N442 , \position1/N441 , \position1/N440 ,
         \position1/N439 , \position1/N438 , \position1/N437 ,
         \position1/N436 , \position1/N435 , \position1/N434 ,
         \position1/N433 , \position1/N432 , \position1/N431 ,
         \position1/N429 , \position1/N428 , \position1/N427 ,
         \position1/N426 , \position1/N425 , \position1/N424 ,
         \position1/N423 , \position1/N422 , \position1/N421 ,
         \position1/N420 , \position1/N419 , \position1/N418 ,
         \position1/N417 , \position1/N416 , \position1/N415 ,
         \position1/N414 , \position1/N413 , \position1/N412 ,
         \position1/N411 , \position1/N410 , \position1/N409 ,
         \position1/N408 , \position1/N407 , \position1/N406 ,
         \position1/N379 , \position1/N378 , \position1/N377 ,
         \position1/N376 , \position1/N375 , \position1/N374 ,
         \position1/N373 , \position1/N372 , \position1/N371 ,
         \position1/N370 , \position1/N369 , \position1/N368 ,
         \position1/N367 , \position1/N366 , \position1/N365 ,
         \position1/N364 , \position1/N363 , \position1/N362 ,
         \position1/N361 , \position1/N360 , \position1/N359 ,
         \position1/N358 , \position1/N357 , \position1/N356 ,
         \position1/N355 , \position1/N354 , \position1/N353 ,
         \position1/N352 , \position1/N351 , \position1/N350 ,
         \position1/N349 , \position1/N348 , \position1/N347 ,
         \position1/N346 , \position1/N345 , \position1/N344 ,
         \position1/N343 , \position1/N342 , \position1/N341 ,
         \position1/N340 , \position1/N339 , \position1/N338 ,
         \position1/N337 , \position1/N336 , \position1/N335 ,
         \position1/N334 , \position1/N333 , \position1/N332 ,
         \position1/N331 , \position1/N304 , \position1/N303 ,
         \position1/N302 , \position1/N301 , \position1/N300 ,
         \position1/N299 , \position1/N298 , \position1/N297 ,
         \position1/N296 , \position1/N295 , \position1/N294 ,
         \position1/N293 , \position1/N292 , \position1/N291 ,
         \position1/N290 , \position1/N289 , \position1/N288 ,
         \position1/N287 , \position1/N286 , \position1/N285 ,
         \position1/N284 , \position1/N283 , \position1/N282 ,
         \position1/N281 , \position1/N280 , \position1/N267 ,
         \position1/N224 , \position1/N223 , \position1/N222 ,
         \position1/N221 , \position1/N220 , \position1/N219 ,
         \position1/N218 , \position1/N217 , \position1/N216 ,
         \position1/N215 , \position1/N214 , \position1/N213 ,
         \position1/N212 , \position1/N211 , \position1/N210 ,
         \position1/N209 , \position1/N208 , \position1/N207 ,
         \position1/N206 , \position1/N194 , \position1/N193 ,
         \position1/N104 , \position1/N103 , \position1/N102 ,
         \position1/N101 , \position1/N100 , \position1/N99 , \position1/N98 ,
         \position1/N97 , \position1/N95 , \position1/N94 , \position1/N93 ,
         \position1/N91 , \position1/N89 , \position1/N88 , \position1/N87 ,
         \position1/N86 , \position1/N85 , \position1/N84 , \position1/N83 ,
         \position1/N82 , \position1/N81 , \position1/r457/carry[2] ,
         \position1/r457/carry[3] , \position1/r457/carry[4] ,
         \position1/r457/carry[5] , \position1/r457/carry[6] ,
         \position1/r457/carry[7] , \position1/r457/carry[8] ,
         \position1/r457/carry[9] , \position1/r457/carry[10] ,
         \position1/r457/carry[11] , \position1/r457/carry[12] ,
         \position1/r457/carry[13] , \position1/r457/carry[14] ,
         \position1/r457/carry[15] , \position1/r457/carry[16] ,
         \position1/r457/carry[17] , \position1/sub_250/carry[2] ,
         \position1/sub_250/carry[3] , \position1/sub_250/carry[4] ,
         \position1/sub_250/carry[5] , \position1/sub_250/carry[6] ,
         \position1/sub_250/carry[7] , \position1/sub_250_3/carry[2] ,
         \position1/sub_250_3/carry[3] , \position1/sub_250_3/carry[4] ,
         \position1/sub_250_3/carry[5] , \position1/sub_250_3/carry[6] ,
         \position1/sub_250_3/carry[7] , \position1/add_250/carry[2] ,
         \position1/add_250/carry[3] , \position1/add_250/carry[4] ,
         \position1/add_250/carry[5] , \position1/add_250/carry[6] ,
         \position1/add_250/carry[7] , \position1/add_250/carry[8] ,
         \position1/add_250_2/carry[2] , \position1/add_250_2/carry[3] ,
         \position1/add_250_2/carry[4] , \position1/add_250_2/carry[5] ,
         \position1/add_250_2/carry[6] , \position1/add_250_2/carry[7] ,
         \position1/add_250_2/carry[8] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[0] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[1] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[2] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[3] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[4] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[5] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[6] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[7] ,
         \position1/dp_cluster_0/mult_add_196_aco/PROD_not[8] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[0] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[1] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[2] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[3] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[4] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[5] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[6] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[7] ,
         \position1/dp_cluster_1/mult_add_197_aco/PROD_not[8] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[0] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[1] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[2] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[3] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[4] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[5] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[6] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[7] ,
         \position1/dp_cluster_4/mult_add_178_aco/PROD_not[8] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[0] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[1] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[2] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[3] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[4] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[5] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[6] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[7] ,
         \position1/dp_cluster_5/mult_add_179_aco/PROD_not[8] ,
         \gensync1/sub_95_2_cf/carry[2] , \gensync1/sub_95_2_cf/carry[3] ,
         \gensync1/sub_95_2_cf/carry[4] , \gensync1/sub_95_2_cf/carry[5] ,
         \gensync1/sub_95_2_cf/carry[6] , \gensync1/sub_95_2_cf/carry[7] ,
         \gensync1/sub_95_2_cf/carry[8] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n491,
         n493, n495, n497, n499, n501, n503, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
  wire   [7:0] \image_process1/bi ;
  wire   [7:0] \image_process1/gi ;
  wire   [7:0] \image_process1/ri ;
  wire   [8:0] \position1/quot_y ;
  wire   [8:0] \position1/quot_x ;
  wire   [1:0] \position1/state ;
  wire   [19:0] \position1/count_img ;
  wire   [24:0] \position1/y_sum ;
  wire   [24:0] \position1/x_sum ;
  wire   [7:0] \position1/gi ;
  wire   [24:1] \position1/r406/carry ;
  wire   [24:1] \position1/r409/carry ;
  wire   [24:1] \position1/r412/carry ;
  wire   [24:1] \position1/r413/carry ;
  wire   [17:2] \position1/r416/carry ;
  wire   [17:1] \position1/r458/carry ;
  wire   [19:2] \position1/add_161/carry ;
  wire   [25:0] \position1/sub_216/carry ;
  wire   [25:0] \position1/sub_216_I2/carry ;
  wire   [25:0] \position1/sub_216_I3/carry ;
  wire   [25:0] \position1/sub_216_I4/carry ;
  wire   [25:0] \position1/sub_216_I5/carry ;
  wire   [25:0] \position1/sub_216_I6/carry ;
  wire   [25:0] \position1/sub_216_I7/carry ;
  wire   [25:0] \position1/sub_216_I8/carry ;
  wire   [25:0] \position1/sub_226/carry ;
  wire   [25:0] \position1/sub_226_I2/carry ;
  wire   [25:0] \position1/sub_226_I3/carry ;
  wire   [25:0] \position1/sub_226_I4/carry ;
  wire   [25:0] \position1/sub_226_I5/carry ;
  wire   [25:0] \position1/sub_226_I6/carry ;
  wire   [25:0] \position1/sub_226_I7/carry ;
  wire   [25:0] \position1/sub_226_I8/carry ;
  wire   [24:1] \position1/dp_cluster_0/add_196_aco/carry ;
  wire   [24:1] \position1/dp_cluster_1/add_197_aco/carry ;
  wire   [24:1] \position1/dp_cluster_2/add_0_root_add_189_3/carry ;
  wire   [24:1] \position1/dp_cluster_3/add_1_root_add_188_3/carry ;
  wire   [24:1] \position1/dp_cluster_3/add_0_root_add_188_3/carry ;
  wire   [24:1] \position1/dp_cluster_4/add_178_aco/carry ;
  wire   [24:1] \position1/dp_cluster_5/add_179_aco/carry ;
  wire   [24:1] \position1/dp_cluster_6/add_1_root_add_171_3/carry ;
  wire   [24:1] \position1/dp_cluster_6/add_0_root_add_171_3/carry ;
  wire   [24:1] \position1/dp_cluster_7/add_1_root_add_170_3/carry ;
  wire   [24:1] \position1/dp_cluster_7/add_0_root_add_170_3/carry ;
  wire   [9:2] \gensync1/add_39/carry ;
  wire   [9:2] \gensync1/add_45/carry ;
  assign cam_x[9] = \*Logic0* ;
  assign cam_x[8] = \position1/dp_cluster_7/N314 ;
  assign cam_y[8] = \position1/dp_cluster_6/N389 ;
  assign cam_y[7] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [8];
  assign cam_y[6] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [7];
  assign cam_y[5] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [6];
  assign cam_y[4] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [5];
  assign cam_y[3] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [4];
  assign cam_y[2] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [3];
  assign cam_y[1] = \position1/dp_cluster_6/add_1_root_add_171_3/carry  [2];

  OAI212 \image_process1/U70  ( .A(n813), .B(\image_process1/n13 ), .C(
        \image_process1/n110 ), .Q(\image_process1/N14 ) );
  OAI212 \image_process1/U68  ( .A(n813), .B(\image_process1/n25 ), .C(
        \image_process1/n110 ), .Q(\image_process1/N16 ) );
  OAI212 \position1/U1019  ( .A(\position1/N1519 ), .B(n97), .C(
        \position1/n1578 ), .Q(\position1/N1573 ) );
  OAI212 \position1/U1017  ( .A(\position1/N1519 ), .B(n91), .C(
        \position1/n1577 ), .Q(\position1/N1547 ) );
  OAI212 \position1/U1015  ( .A(n518), .B(n90), .C(\position1/n1576 ), .Q(
        \position1/N1548 ) );
  OAI212 \position1/U1013  ( .A(n520), .B(n95), .C(\position1/n1575 ), .Q(
        \position1/N1549 ) );
  OAI212 \position1/U1011  ( .A(n520), .B(n89), .C(\position1/n1574 ), .Q(
        \position1/N1550 ) );
  OAI212 \position1/U1009  ( .A(n520), .B(n88), .C(\position1/n1573 ), .Q(
        \position1/N1551 ) );
  OAI212 \position1/U1007  ( .A(n520), .B(n87), .C(\position1/n1572 ), .Q(
        \position1/N1552 ) );
  OAI212 \position1/U1005  ( .A(n520), .B(n94), .C(\position1/n1571 ), .Q(
        \position1/N1553 ) );
  OAI212 \position1/U1003  ( .A(n520), .B(n49), .C(\position1/n1570 ), .Q(
        \position1/N1554 ) );
  OAI212 \position1/U1001  ( .A(n520), .B(n51), .C(\position1/n1569 ), .Q(
        \position1/N1555 ) );
  OAI212 \position1/U999  ( .A(n520), .B(n69), .C(\position1/n1568 ), .Q(
        \position1/N1556 ) );
  OAI212 \position1/U997  ( .A(n520), .B(n65), .C(\position1/n1567 ), .Q(
        \position1/N1557 ) );
  OAI212 \position1/U995  ( .A(n520), .B(n81), .C(\position1/n1566 ), .Q(
        \position1/N1558 ) );
  OAI212 \position1/U993  ( .A(n520), .B(n64), .C(\position1/n1565 ), .Q(
        \position1/N1559 ) );
  OAI212 \position1/U991  ( .A(n520), .B(n80), .C(\position1/n1564 ), .Q(
        \position1/N1560 ) );
  OAI212 \position1/U989  ( .A(n520), .B(n63), .C(\position1/n1563 ), .Q(
        \position1/N1561 ) );
  OAI212 \position1/U987  ( .A(n520), .B(n79), .C(\position1/n1562 ), .Q(
        \position1/N1562 ) );
  OAI212 \position1/U985  ( .A(n520), .B(n62), .C(\position1/n1561 ), .Q(
        \position1/N1563 ) );
  OAI212 \position1/U983  ( .A(n520), .B(n78), .C(\position1/n1560 ), .Q(
        \position1/N1564 ) );
  OAI212 \position1/U981  ( .A(n519), .B(n61), .C(\position1/n1559 ), .Q(
        \position1/N1565 ) );
  OAI212 \position1/U979  ( .A(n519), .B(n77), .C(\position1/n1558 ), .Q(
        \position1/N1566 ) );
  OAI212 \position1/U977  ( .A(n518), .B(n60), .C(\position1/n1557 ), .Q(
        \position1/N1567 ) );
  OAI212 \position1/U975  ( .A(\position1/N1519 ), .B(n76), .C(
        \position1/n1556 ), .Q(\position1/N1568 ) );
  OAI212 \position1/U973  ( .A(\position1/N1519 ), .B(n59), .C(
        \position1/n1555 ), .Q(\position1/N1569 ) );
  OAI212 \position1/U971  ( .A(\position1/N1519 ), .B(n99), .C(
        \position1/n1554 ), .Q(\position1/N1570 ) );
  OAI222 \position1/U945  ( .A(n528), .B(\position1/n1553 ), .C(n526), .D(
        \position1/n1553 ), .Q(\position1/N1677 ) );
  OAI222 \position1/U944  ( .A(n529), .B(\position1/n1552 ), .C(n526), .D(
        \position1/n1552 ), .Q(\position1/N1651 ) );
  OAI222 \position1/U943  ( .A(n529), .B(\position1/n1551 ), .C(n526), .D(
        \position1/n1551 ), .Q(\position1/N1652 ) );
  OAI222 \position1/U942  ( .A(n529), .B(\position1/n1550 ), .C(n526), .D(
        \position1/n1550 ), .Q(\position1/N1653 ) );
  OAI222 \position1/U941  ( .A(n529), .B(\position1/n1549 ), .C(n526), .D(
        \position1/n1549 ), .Q(\position1/N1654 ) );
  OAI222 \position1/U940  ( .A(n529), .B(\position1/n1548 ), .C(n526), .D(
        \position1/n1548 ), .Q(\position1/N1655 ) );
  OAI222 \position1/U939  ( .A(n529), .B(n104), .C(n526), .D(\position1/n1547 ), .Q(\position1/N1656 ) );
  OAI222 \position1/U938  ( .A(n529), .B(n1297), .C(n526), .D(
        \position1/n1546 ), .Q(\position1/N1657 ) );
  OAI222 \position1/U937  ( .A(n529), .B(n1294), .C(n526), .D(
        \position1/n1545 ), .Q(\position1/N1658 ) );
  OAI222 \position1/U936  ( .A(n529), .B(n1292), .C(n526), .D(
        \position1/n1544 ), .Q(\position1/N1659 ) );
  OAI222 \position1/U935  ( .A(n529), .B(n1289), .C(n526), .D(
        \position1/n1543 ), .Q(\position1/N1660 ) );
  OAI222 \position1/U934  ( .A(n530), .B(n1287), .C(n526), .D(
        \position1/n1542 ), .Q(\position1/N1661 ) );
  OAI222 \position1/U933  ( .A(n530), .B(n1285), .C(n526), .D(
        \position1/n1541 ), .Q(\position1/N1662 ) );
  OAI222 \position1/U932  ( .A(n530), .B(n1283), .C(n527), .D(
        \position1/n1540 ), .Q(\position1/N1663 ) );
  OAI222 \position1/U931  ( .A(n530), .B(n1281), .C(n527), .D(
        \position1/n1539 ), .Q(\position1/N1664 ) );
  OAI222 \position1/U930  ( .A(n528), .B(n1279), .C(n527), .D(
        \position1/n1538 ), .Q(\position1/N1665 ) );
  OAI222 \position1/U929  ( .A(n530), .B(n1277), .C(n527), .D(
        \position1/n1537 ), .Q(\position1/N1666 ) );
  OAI222 \position1/U928  ( .A(n528), .B(n1275), .C(n527), .D(
        \position1/n1536 ), .Q(\position1/N1667 ) );
  OAI222 \position1/U927  ( .A(n530), .B(n1273), .C(n527), .D(
        \position1/n1535 ), .Q(\position1/N1668 ) );
  OAI222 \position1/U926  ( .A(n530), .B(n1271), .C(n527), .D(
        \position1/n1534 ), .Q(\position1/N1669 ) );
  OAI222 \position1/U925  ( .A(n530), .B(n1269), .C(n527), .D(
        \position1/n1533 ), .Q(\position1/N1670 ) );
  OAI222 \position1/U924  ( .A(n528), .B(n1248), .C(n527), .D(
        \position1/n1532 ), .Q(\position1/N1671 ) );
  OAI222 \position1/U923  ( .A(n528), .B(n1246), .C(n527), .D(
        \position1/n1531 ), .Q(\position1/N1672 ) );
  OAI222 \position1/U922  ( .A(n528), .B(n1245), .C(n527), .D(
        \position1/n1530 ), .Q(\position1/N1673 ) );
  OAI222 \position1/U921  ( .A(n528), .B(n106), .C(n527), .D(\position1/n1529 ), .Q(\position1/N1674 ) );
  OAI212 \position1/U799  ( .A(\position1/state [1]), .B(\position1/state [0]), 
        .C(n486), .Q(\position1/N2353 ) );
  OAI212 \position1/U783  ( .A(\position1/n1395 ), .B(\position1/n1396 ), .C(
        n851), .Q(\position1/n1390 ) );
  OAI222 \position1/U773  ( .A(n1358), .B(n652), .C(\position1/n1141 ), .D(
        \position1/n1064 ), .Q(\position1/N193 ) );
  OAI212 \position1/U764  ( .A(\position1/N1936 ), .B(n96), .C(
        \position1/n1382 ), .Q(\position1/N1990 ) );
  OAI212 \position1/U762  ( .A(\position1/N1936 ), .B(n86), .C(
        \position1/n1381 ), .Q(\position1/N1964 ) );
  OAI212 \position1/U760  ( .A(n552), .B(n85), .C(\position1/n1380 ), .Q(
        \position1/N1965 ) );
  OAI212 \position1/U758  ( .A(n554), .B(n93), .C(\position1/n1379 ), .Q(
        \position1/N1966 ) );
  OAI212 \position1/U756  ( .A(n554), .B(n84), .C(\position1/n1378 ), .Q(
        \position1/N1967 ) );
  OAI212 \position1/U754  ( .A(n554), .B(n83), .C(\position1/n1377 ), .Q(
        \position1/N1968 ) );
  OAI212 \position1/U752  ( .A(n554), .B(n82), .C(\position1/n1376 ), .Q(
        \position1/N1969 ) );
  OAI212 \position1/U750  ( .A(n554), .B(n92), .C(\position1/n1375 ), .Q(
        \position1/N1970 ) );
  OAI212 \position1/U748  ( .A(n554), .B(n48), .C(\position1/n1374 ), .Q(
        \position1/N1971 ) );
  OAI212 \position1/U746  ( .A(n554), .B(n50), .C(\position1/n1373 ), .Q(
        \position1/N1972 ) );
  OAI212 \position1/U744  ( .A(n554), .B(n68), .C(\position1/n1372 ), .Q(
        \position1/N1973 ) );
  OAI212 \position1/U742  ( .A(n554), .B(n58), .C(\position1/n1371 ), .Q(
        \position1/N1974 ) );
  OAI212 \position1/U740  ( .A(n554), .B(n75), .C(\position1/n1370 ), .Q(
        \position1/N1975 ) );
  OAI212 \position1/U738  ( .A(n554), .B(n57), .C(\position1/n1369 ), .Q(
        \position1/N1976 ) );
  OAI212 \position1/U736  ( .A(n554), .B(n74), .C(\position1/n1368 ), .Q(
        \position1/N1977 ) );
  OAI212 \position1/U734  ( .A(n554), .B(n56), .C(\position1/n1367 ), .Q(
        \position1/N1978 ) );
  OAI212 \position1/U732  ( .A(n554), .B(n73), .C(\position1/n1366 ), .Q(
        \position1/N1979 ) );
  OAI212 \position1/U730  ( .A(n554), .B(n55), .C(\position1/n1365 ), .Q(
        \position1/N1980 ) );
  OAI212 \position1/U728  ( .A(n554), .B(n72), .C(\position1/n1364 ), .Q(
        \position1/N1981 ) );
  OAI212 \position1/U726  ( .A(n553), .B(n54), .C(\position1/n1363 ), .Q(
        \position1/N1982 ) );
  OAI212 \position1/U724  ( .A(n553), .B(n71), .C(\position1/n1362 ), .Q(
        \position1/N1983 ) );
  OAI212 \position1/U722  ( .A(n552), .B(n53), .C(\position1/n1361 ), .Q(
        \position1/N1984 ) );
  OAI212 \position1/U720  ( .A(\position1/N1936 ), .B(n70), .C(
        \position1/n1360 ), .Q(\position1/N1985 ) );
  OAI212 \position1/U718  ( .A(\position1/N1936 ), .B(n52), .C(
        \position1/n1359 ), .Q(\position1/N1986 ) );
  OAI212 \position1/U716  ( .A(\position1/N1936 ), .B(n98), .C(
        \position1/n1358 ), .Q(\position1/N1987 ) );
  OAI222 \position1/U690  ( .A(n562), .B(\position1/n1357 ), .C(n560), .D(
        \position1/n1357 ), .Q(\position1/N2094 ) );
  OAI222 \position1/U689  ( .A(n563), .B(\position1/n1356 ), .C(n560), .D(
        \position1/n1356 ), .Q(\position1/N2068 ) );
  OAI222 \position1/U688  ( .A(n563), .B(\position1/n1355 ), .C(n560), .D(
        \position1/n1355 ), .Q(\position1/N2069 ) );
  OAI222 \position1/U687  ( .A(n563), .B(\position1/n1354 ), .C(n560), .D(
        \position1/n1354 ), .Q(\position1/N2070 ) );
  OAI222 \position1/U686  ( .A(n563), .B(\position1/n1353 ), .C(n560), .D(
        \position1/n1353 ), .Q(\position1/N2071 ) );
  OAI222 \position1/U685  ( .A(n563), .B(\position1/n1352 ), .C(n560), .D(
        \position1/n1352 ), .Q(\position1/N2072 ) );
  OAI222 \position1/U684  ( .A(n563), .B(n105), .C(n560), .D(\position1/n1351 ), .Q(\position1/N2073 ) );
  OAI222 \position1/U683  ( .A(n563), .B(n1078), .C(n560), .D(
        \position1/n1350 ), .Q(\position1/N2074 ) );
  OAI222 \position1/U682  ( .A(n563), .B(n1075), .C(n560), .D(
        \position1/n1349 ), .Q(\position1/N2075 ) );
  OAI222 \position1/U681  ( .A(n563), .B(n1073), .C(n560), .D(
        \position1/n1348 ), .Q(\position1/N2076 ) );
  OAI222 \position1/U680  ( .A(n563), .B(n1070), .C(n560), .D(
        \position1/n1347 ), .Q(\position1/N2077 ) );
  OAI222 \position1/U679  ( .A(n564), .B(n1068), .C(n560), .D(
        \position1/n1346 ), .Q(\position1/N2078 ) );
  OAI222 \position1/U678  ( .A(n564), .B(n1066), .C(n560), .D(
        \position1/n1345 ), .Q(\position1/N2079 ) );
  OAI222 \position1/U677  ( .A(n564), .B(n1064), .C(n561), .D(
        \position1/n1344 ), .Q(\position1/N2080 ) );
  OAI222 \position1/U676  ( .A(n564), .B(n1062), .C(n561), .D(
        \position1/n1343 ), .Q(\position1/N2081 ) );
  OAI222 \position1/U675  ( .A(n562), .B(n1060), .C(n561), .D(
        \position1/n1342 ), .Q(\position1/N2082 ) );
  OAI222 \position1/U674  ( .A(n564), .B(n1058), .C(n561), .D(
        \position1/n1341 ), .Q(\position1/N2083 ) );
  OAI222 \position1/U673  ( .A(n562), .B(n1056), .C(n561), .D(
        \position1/n1340 ), .Q(\position1/N2084 ) );
  OAI222 \position1/U672  ( .A(n564), .B(n1054), .C(n561), .D(
        \position1/n1339 ), .Q(\position1/N2085 ) );
  OAI222 \position1/U671  ( .A(n564), .B(n1052), .C(n561), .D(
        \position1/n1338 ), .Q(\position1/N2086 ) );
  OAI222 \position1/U670  ( .A(n564), .B(n1050), .C(n561), .D(
        \position1/n1337 ), .Q(\position1/N2087 ) );
  OAI222 \position1/U669  ( .A(n562), .B(n1029), .C(n561), .D(
        \position1/n1336 ), .Q(\position1/N2088 ) );
  OAI222 \position1/U668  ( .A(n562), .B(n1027), .C(n561), .D(
        \position1/n1335 ), .Q(\position1/N2089 ) );
  OAI222 \position1/U667  ( .A(n562), .B(n1026), .C(n561), .D(
        \position1/n1334 ), .Q(\position1/N2090 ) );
  OAI222 \position1/U666  ( .A(n562), .B(n107), .C(n561), .D(\position1/n1333 ), .Q(\position1/N2091 ) );
  OAI212 \position1/U487  ( .A(n654), .B(\position1/n362 ), .C(n712), .Q(
        \position1/N89 ) );
  OAI212 \position1/U485  ( .A(n654), .B(\position1/n360 ), .C(n712), .Q(
        \position1/N91 ) );
  OAI212 \position1/U483  ( .A(n653), .B(\position1/n358 ), .C(n712), .Q(
        \position1/N93 ) );
  OAI212 \position1/U482  ( .A(n652), .B(\position1/n357 ), .C(n712), .Q(
        \position1/N94 ) );
  OAI212 \position1/U481  ( .A(n652), .B(\position1/n356 ), .C(n712), .Q(
        \position1/N95 ) );
  OAI222 \position1/U447  ( .A(\position1/n1063 ), .B(\position1/n1151 ), .C(
        \position1/n1141 ), .D(\position1/n1145 ), .Q(\position1/n1072 ) );
  OAI222 \position1/U445  ( .A(\position1/n1149 ), .B(\position1/n1062 ), .C(
        \position1/n1146 ), .D(\position1/n1141 ), .Q(\position1/n1060 ) );
  OAI222 \position1/U438  ( .A(\position1/n1062 ), .B(\position1/n1065 ), .C(
        \position1/n1141 ), .D(\position1/n1058 ), .Q(\position1/n1071 ) );
  ADD32 \position1/r406/U1_1  ( .A(\position1/x_sum [1]), .B(cam_x[1]), .CI(
        \position1/r406/carry [1]), .CO(\position1/r406/carry [2]), .S(
        \position1/N281 ) );
  ADD32 \position1/r406/U1_2  ( .A(\position1/x_sum [2]), .B(cam_x[2]), .CI(
        \position1/r406/carry [2]), .CO(\position1/r406/carry [3]), .S(
        \position1/N282 ) );
  ADD32 \position1/r406/U1_3  ( .A(\position1/x_sum [3]), .B(cam_x[3]), .CI(
        \position1/r406/carry [3]), .CO(\position1/r406/carry [4]), .S(
        \position1/N283 ) );
  ADD32 \position1/r406/U1_4  ( .A(\position1/x_sum [4]), .B(cam_x[4]), .CI(
        \position1/r406/carry [4]), .CO(\position1/r406/carry [5]), .S(
        \position1/N284 ) );
  ADD32 \position1/r406/U1_5  ( .A(\position1/x_sum [5]), .B(cam_x[5]), .CI(
        \position1/r406/carry [5]), .CO(\position1/r406/carry [6]), .S(
        \position1/N285 ) );
  ADD32 \position1/r406/U1_6  ( .A(\position1/x_sum [6]), .B(cam_x[6]), .CI(
        \position1/r406/carry [6]), .CO(\position1/r406/carry [7]), .S(
        \position1/N286 ) );
  ADD32 \position1/r406/U1_7  ( .A(\position1/x_sum [7]), .B(cam_x[7]), .CI(
        \position1/r406/carry [7]), .CO(\position1/r406/carry [8]), .S(
        \position1/N287 ) );
  ADD32 \position1/r406/U1_8  ( .A(\position1/x_sum [8]), .B(
        \position1/dp_cluster_7/N314 ), .CI(\position1/r406/carry [8]), .CO(
        \position1/r406/carry [9]), .S(\position1/N288 ) );
  ADD32 \position1/r409/U1_1  ( .A(\position1/y_sum [1]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .CI(
        \position1/r409/carry [1]), .CO(\position1/r409/carry [2]), .S(
        \position1/N356 ) );
  ADD32 \position1/r409/U1_2  ( .A(\position1/y_sum [2]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .CI(
        \position1/r409/carry [2]), .CO(\position1/r409/carry [3]), .S(
        \position1/N357 ) );
  ADD32 \position1/r409/U1_3  ( .A(\position1/y_sum [3]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), .CI(
        \position1/r409/carry [3]), .CO(\position1/r409/carry [4]), .S(
        \position1/N358 ) );
  ADD32 \position1/r409/U1_4  ( .A(\position1/y_sum [4]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .CI(
        \position1/r409/carry [4]), .CO(\position1/r409/carry [5]), .S(
        \position1/N359 ) );
  ADD32 \position1/r409/U1_5  ( .A(\position1/y_sum [5]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .CI(
        \position1/r409/carry [5]), .CO(\position1/r409/carry [6]), .S(
        \position1/N360 ) );
  ADD32 \position1/r409/U1_6  ( .A(\position1/y_sum [6]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .CI(
        \position1/r409/carry [6]), .CO(\position1/r409/carry [7]), .S(
        \position1/N361 ) );
  ADD32 \position1/r409/U1_7  ( .A(\position1/y_sum [7]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .CI(
        \position1/r409/carry [7]), .CO(\position1/r409/carry [8]), .S(
        \position1/N362 ) );
  ADD32 \position1/r409/U1_8  ( .A(\position1/y_sum [8]), .B(
        \position1/dp_cluster_6/N389 ), .CI(\position1/r409/carry [8]), .CO(
        \position1/r409/carry [9]), .S(\position1/N363 ) );
  ADD32 \position1/r412/U1_1  ( .A(n501), .B(\position1/N281 ), .CI(
        \position1/r412/carry [1]), .CO(\position1/r412/carry [2]), .S(
        \position1/N486 ) );
  ADD32 \position1/r412/U1_2  ( .A(n499), .B(\position1/N282 ), .CI(
        \position1/r412/carry [2]), .CO(\position1/r412/carry [3]), .S(
        \position1/N487 ) );
  ADD32 \position1/r412/U1_3  ( .A(n497), .B(\position1/N283 ), .CI(
        \position1/r412/carry [3]), .CO(\position1/r412/carry [4]), .S(
        \position1/N488 ) );
  ADD32 \position1/r412/U1_4  ( .A(n495), .B(\position1/N284 ), .CI(
        \position1/r412/carry [4]), .CO(\position1/r412/carry [5]), .S(
        \position1/N489 ) );
  ADD32 \position1/r412/U1_5  ( .A(n493), .B(\position1/N285 ), .CI(
        \position1/r412/carry [5]), .CO(\position1/r412/carry [6]), .S(
        \position1/N490 ) );
  ADD32 \position1/r412/U1_6  ( .A(n491), .B(\position1/N286 ), .CI(
        \position1/r412/carry [6]), .CO(\position1/r412/carry [7]), .S(
        \position1/N491 ) );
  ADD32 \position1/r412/U1_7  ( .A(n489), .B(\position1/N287 ), .CI(
        \position1/r412/carry [7]), .CO(\position1/r412/carry [8]), .S(
        \position1/N492 ) );
  ADD32 \position1/r412/U1_8  ( .A(\position1/dp_cluster_7/N314 ), .B(
        \position1/N288 ), .CI(\position1/r412/carry [8]), .CO(
        \position1/r412/carry [9]), .S(\position1/N493 ) );
  ADD32 \position1/r413/U1_1  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .B(
        \position1/N356 ), .CI(\position1/r413/carry [1]), .CO(
        \position1/r413/carry [2]), .S(\position1/N536 ) );
  ADD32 \position1/r413/U1_2  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .B(
        \position1/N357 ), .CI(\position1/r413/carry [2]), .CO(
        \position1/r413/carry [3]), .S(\position1/N537 ) );
  ADD32 \position1/r413/U1_3  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), .B(
        \position1/N358 ), .CI(\position1/r413/carry [3]), .CO(
        \position1/r413/carry [4]), .S(\position1/N538 ) );
  ADD32 \position1/r413/U1_4  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .B(
        \position1/N359 ), .CI(\position1/r413/carry [4]), .CO(
        \position1/r413/carry [5]), .S(\position1/N539 ) );
  ADD32 \position1/r413/U1_5  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .B(
        \position1/N360 ), .CI(\position1/r413/carry [5]), .CO(
        \position1/r413/carry [6]), .S(\position1/N540 ) );
  ADD32 \position1/r413/U1_6  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .B(
        \position1/N361 ), .CI(\position1/r413/carry [6]), .CO(
        \position1/r413/carry [7]), .S(\position1/N541 ) );
  ADD32 \position1/r413/U1_7  ( .A(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .B(
        \position1/N362 ), .CI(\position1/r413/carry [7]), .CO(
        \position1/r413/carry [8]), .S(\position1/N542 ) );
  ADD32 \position1/r413/U1_8  ( .A(\position1/dp_cluster_6/N389 ), .B(
        \position1/N363 ), .CI(\position1/r413/carry [8]), .CO(
        \position1/r413/carry [9]), .S(\position1/N543 ) );
  ADD22 \position1/r416/U1_1_1  ( .A(n631), .B(n514), .CO(
        \position1/r416/carry [2]), .S(\position1/N590 ) );
  ADD22 \position1/r416/U1_1_2  ( .A(n627), .B(\position1/r416/carry [2]), 
        .CO(\position1/r416/carry [3]), .S(\position1/N591 ) );
  ADD22 \position1/r416/U1_1_3  ( .A(n623), .B(\position1/r416/carry [3]), 
        .CO(\position1/r416/carry [4]), .S(\position1/N592 ) );
  ADD22 \position1/r416/U1_1_4  ( .A(n468), .B(\position1/r416/carry [4]), 
        .CO(\position1/r416/carry [5]), .S(\position1/N593 ) );
  ADD22 \position1/r416/U1_1_5  ( .A(n620), .B(\position1/r416/carry [5]), 
        .CO(\position1/r416/carry [6]), .S(\position1/N594 ) );
  ADD22 \position1/r416/U1_1_6  ( .A(n469), .B(\position1/r416/carry [6]), 
        .CO(\position1/r416/carry [7]), .S(\position1/N595 ) );
  ADD22 \position1/r416/U1_1_7  ( .A(n615), .B(\position1/r416/carry [7]), 
        .CO(\position1/r416/carry [8]), .S(\position1/N596 ) );
  ADD22 \position1/r416/U1_1_8  ( .A(n471), .B(\position1/r416/carry [8]), 
        .CO(\position1/r416/carry [9]), .S(\position1/N597 ) );
  ADD22 \position1/r416/U1_1_9  ( .A(n608), .B(\position1/r416/carry [9]), 
        .CO(\position1/r416/carry [10]), .S(\position1/N598 ) );
  ADD22 \position1/r416/U1_1_10  ( .A(n473), .B(\position1/r416/carry [10]), 
        .CO(\position1/r416/carry [11]), .S(\position1/N599 ) );
  ADD22 \position1/r416/U1_1_11  ( .A(n605), .B(\position1/r416/carry [11]), 
        .CO(\position1/r416/carry [12]), .S(\position1/N600 ) );
  ADD22 \position1/r416/U1_1_12  ( .A(n474), .B(\position1/r416/carry [12]), 
        .CO(\position1/r416/carry [13]), .S(\position1/N601 ) );
  ADD22 \position1/r416/U1_1_13  ( .A(n601), .B(\position1/r416/carry [13]), 
        .CO(\position1/r416/carry [14]), .S(\position1/N602 ) );
  ADD22 \position1/r416/U1_1_14  ( .A(n475), .B(\position1/r416/carry [14]), 
        .CO(\position1/r416/carry [15]), .S(\position1/N603 ) );
  ADD22 \position1/r416/U1_1_15  ( .A(n597), .B(\position1/r416/carry [15]), 
        .CO(\position1/r416/carry [16]), .S(\position1/N604 ) );
  ADD22 \position1/r416/U1_1_16  ( .A(n594), .B(\position1/r416/carry [16]), 
        .CO(\position1/r416/carry [17]), .S(\position1/N605 ) );
  ADD22 \position1/add_161/U1_1_1  ( .A(\position1/count_img [1]), .B(
        \position1/count_img [0]), .CO(\position1/add_161/carry [2]), .S(
        \position1/N206 ) );
  ADD22 \position1/add_161/U1_1_2  ( .A(\position1/count_img [2]), .B(
        \position1/add_161/carry [2]), .CO(\position1/add_161/carry [3]), .S(
        \position1/N207 ) );
  ADD22 \position1/add_161/U1_1_3  ( .A(\position1/count_img [3]), .B(
        \position1/add_161/carry [3]), .CO(\position1/add_161/carry [4]), .S(
        \position1/N208 ) );
  ADD22 \position1/add_161/U1_1_4  ( .A(\position1/count_img [4]), .B(
        \position1/add_161/carry [4]), .CO(\position1/add_161/carry [5]), .S(
        \position1/N209 ) );
  ADD22 \position1/add_161/U1_1_5  ( .A(\position1/count_img [5]), .B(
        \position1/add_161/carry [5]), .CO(\position1/add_161/carry [6]), .S(
        \position1/N210 ) );
  ADD22 \position1/add_161/U1_1_6  ( .A(\position1/count_img [6]), .B(
        \position1/add_161/carry [6]), .CO(\position1/add_161/carry [7]), .S(
        \position1/N211 ) );
  ADD22 \position1/add_161/U1_1_7  ( .A(\position1/count_img [7]), .B(
        \position1/add_161/carry [7]), .CO(\position1/add_161/carry [8]), .S(
        \position1/N212 ) );
  ADD22 \position1/add_161/U1_1_8  ( .A(\position1/count_img [8]), .B(
        \position1/add_161/carry [8]), .CO(\position1/add_161/carry [9]), .S(
        \position1/N213 ) );
  ADD22 \position1/add_161/U1_1_9  ( .A(\position1/count_img [9]), .B(
        \position1/add_161/carry [9]), .CO(\position1/add_161/carry [10]), .S(
        \position1/N214 ) );
  ADD22 \position1/add_161/U1_1_10  ( .A(\position1/count_img [10]), .B(
        \position1/add_161/carry [10]), .CO(\position1/add_161/carry [11]), 
        .S(\position1/N215 ) );
  ADD22 \position1/add_161/U1_1_11  ( .A(\position1/count_img [11]), .B(
        \position1/add_161/carry [11]), .CO(\position1/add_161/carry [12]), 
        .S(\position1/N216 ) );
  ADD22 \position1/add_161/U1_1_12  ( .A(\position1/count_img [12]), .B(
        \position1/add_161/carry [12]), .CO(\position1/add_161/carry [13]), 
        .S(\position1/N217 ) );
  ADD22 \position1/add_161/U1_1_13  ( .A(\position1/count_img [13]), .B(
        \position1/add_161/carry [13]), .CO(\position1/add_161/carry [14]), 
        .S(\position1/N218 ) );
  ADD22 \position1/add_161/U1_1_14  ( .A(\position1/count_img [14]), .B(
        \position1/add_161/carry [14]), .CO(\position1/add_161/carry [15]), 
        .S(\position1/N219 ) );
  ADD22 \position1/add_161/U1_1_15  ( .A(\position1/count_img [15]), .B(
        \position1/add_161/carry [15]), .CO(\position1/add_161/carry [16]), 
        .S(\position1/N220 ) );
  ADD22 \position1/add_161/U1_1_16  ( .A(\position1/count_img [16]), .B(
        \position1/add_161/carry [16]), .CO(\position1/add_161/carry [17]), 
        .S(\position1/N221 ) );
  ADD22 \position1/add_161/U1_1_17  ( .A(\position1/count_img [17]), .B(
        \position1/add_161/carry [17]), .CO(\position1/add_161/carry [18]), 
        .S(\position1/N222 ) );
  ADD22 \position1/add_161/U1_1_18  ( .A(\position1/count_img [18]), .B(
        \position1/add_161/carry [18]), .CO(\position1/add_161/carry [19]), 
        .S(\position1/N223 ) );
  ADD32 \position1/sub_216/U2_9  ( .A(\position1/x_sum [9]), .B(n628), .CI(
        \position1/sub_216/carry [9]), .CO(\position1/sub_216/carry [10]), .S(
        \position1/N1530 ) );
  ADD32 \position1/sub_216/U2_10  ( .A(\position1/x_sum [10]), .B(n66), .CI(
        \position1/sub_216/carry [10]), .CO(\position1/sub_216/carry [11]), 
        .S(\position1/N1531 ) );
  ADD32 \position1/sub_216/U2_11  ( .A(\position1/x_sum [11]), .B(n274), .CI(
        \position1/sub_216/carry [11]), .CO(\position1/sub_216/carry [12]), 
        .S(\position1/N1532 ) );
  ADD32 \position1/sub_216/U2_12  ( .A(\position1/x_sum [12]), .B(n41), .CI(
        \position1/sub_216/carry [12]), .CO(\position1/sub_216/carry [13]), 
        .S(\position1/N1533 ) );
  ADD32 \position1/sub_216/U2_13  ( .A(\position1/x_sum [13]), .B(n278), .CI(
        \position1/sub_216/carry [13]), .CO(\position1/sub_216/carry [14]), 
        .S(\position1/N1534 ) );
  ADD32 \position1/sub_216/U2_14  ( .A(\position1/x_sum [14]), .B(n280), .CI(
        \position1/sub_216/carry [14]), .CO(\position1/sub_216/carry [15]), 
        .S(\position1/N1535 ) );
  ADD32 \position1/sub_216/U2_15  ( .A(\position1/x_sum [15]), .B(n282), .CI(
        \position1/sub_216/carry [15]), .CO(\position1/sub_216/carry [16]), 
        .S(\position1/N1536 ) );
  ADD32 \position1/sub_216/U2_16  ( .A(\position1/x_sum [16]), .B(n40), .CI(
        \position1/sub_216/carry [16]), .CO(\position1/sub_216/carry [17]), 
        .S(\position1/N1537 ) );
  ADD32 \position1/sub_216/U2_17  ( .A(\position1/x_sum [17]), .B(n286), .CI(
        \position1/sub_216/carry [17]), .CO(\position1/sub_216/carry [18]), 
        .S(\position1/N1538 ) );
  ADD32 \position1/sub_216/U2_18  ( .A(\position1/x_sum [18]), .B(n46), .CI(
        \position1/sub_216/carry [18]), .CO(\position1/sub_216/carry [19]), 
        .S(\position1/N1539 ) );
  ADD32 \position1/sub_216/U2_19  ( .A(\position1/x_sum [19]), .B(n290), .CI(
        \position1/sub_216/carry [19]), .CO(\position1/sub_216/carry [20]), 
        .S(\position1/N1540 ) );
  ADD32 \position1/sub_216/U2_20  ( .A(\position1/x_sum [20]), .B(n43), .CI(
        \position1/sub_216/carry [20]), .CO(\position1/sub_216/carry [21]), 
        .S(\position1/N1541 ) );
  ADD32 \position1/sub_216/U2_21  ( .A(\position1/x_sum [21]), .B(n294), .CI(
        \position1/sub_216/carry [21]), .CO(\position1/sub_216/carry [22]), 
        .S(\position1/N1542 ) );
  ADD32 \position1/sub_216/U2_22  ( .A(\position1/x_sum [22]), .B(n42), .CI(
        \position1/sub_216/carry [22]), .CO(\position1/sub_216/carry [23]), 
        .S(\position1/N1543 ) );
  ADD32 \position1/sub_216/U2_23  ( .A(\position1/x_sum [23]), .B(n298), .CI(
        \position1/sub_216/carry [23]), .CO(\position1/sub_216/carry [24]), 
        .S(\position1/N1544 ) );
  ADD32 \position1/sub_216_I2/U2_8  ( .A(\position1/N1554 ), .B(n36), .CI(
        \position1/sub_216_I2/carry [8]), .CO(\position1/sub_216_I2/carry [9]), 
        .S(\position1/N1581 ) );
  ADD32 \position1/sub_216_I2/U2_9  ( .A(\position1/N1555 ), .B(n272), .CI(
        \position1/sub_216_I2/carry [9]), .CO(\position1/sub_216_I2/carry [10]), .S(\position1/N1582 ) );
  ADD32 \position1/sub_216_I2/U2_10  ( .A(\position1/N1556 ), .B(n274), .CI(
        \position1/sub_216_I2/carry [10]), .CO(
        \position1/sub_216_I2/carry [11]), .S(\position1/N1583 ) );
  ADD32 \position1/sub_216_I2/U2_11  ( .A(\position1/N1557 ), .B(n276), .CI(
        \position1/sub_216_I2/carry [11]), .CO(
        \position1/sub_216_I2/carry [12]), .S(\position1/N1584 ) );
  ADD32 \position1/sub_216_I2/U2_12  ( .A(\position1/N1558 ), .B(n278), .CI(
        \position1/sub_216_I2/carry [12]), .CO(
        \position1/sub_216_I2/carry [13]), .S(\position1/N1585 ) );
  ADD32 \position1/sub_216_I2/U2_13  ( .A(\position1/N1559 ), .B(n280), .CI(
        \position1/sub_216_I2/carry [13]), .CO(
        \position1/sub_216_I2/carry [14]), .S(\position1/N1586 ) );
  ADD32 \position1/sub_216_I2/U2_14  ( .A(\position1/N1560 ), .B(n282), .CI(
        \position1/sub_216_I2/carry [14]), .CO(
        \position1/sub_216_I2/carry [15]), .S(\position1/N1587 ) );
  ADD32 \position1/sub_216_I2/U2_15  ( .A(\position1/N1561 ), .B(n256), .CI(
        \position1/sub_216_I2/carry [15]), .CO(
        \position1/sub_216_I2/carry [16]), .S(\position1/N1588 ) );
  ADD32 \position1/sub_216_I2/U2_16  ( .A(\position1/N1562 ), .B(n35), .CI(
        \position1/sub_216_I2/carry [16]), .CO(
        \position1/sub_216_I2/carry [17]), .S(\position1/N1589 ) );
  ADD32 \position1/sub_216_I2/U2_17  ( .A(\position1/N1563 ), .B(n288), .CI(
        \position1/sub_216_I2/carry [17]), .CO(
        \position1/sub_216_I2/carry [18]), .S(\position1/N1590 ) );
  ADD32 \position1/sub_216_I2/U2_18  ( .A(\position1/N1564 ), .B(n290), .CI(
        \position1/sub_216_I2/carry [18]), .CO(
        \position1/sub_216_I2/carry [19]), .S(\position1/N1591 ) );
  ADD32 \position1/sub_216_I2/U2_19  ( .A(\position1/N1565 ), .B(n263), .CI(
        \position1/sub_216_I2/carry [19]), .CO(
        \position1/sub_216_I2/carry [20]), .S(\position1/N1592 ) );
  ADD32 \position1/sub_216_I2/U2_20  ( .A(\position1/N1566 ), .B(n294), .CI(
        \position1/sub_216_I2/carry [20]), .CO(
        \position1/sub_216_I2/carry [21]), .S(\position1/N1593 ) );
  ADD32 \position1/sub_216_I2/U2_21  ( .A(\position1/N1567 ), .B(n296), .CI(
        \position1/sub_216_I2/carry [21]), .CO(
        \position1/sub_216_I2/carry [22]), .S(\position1/N1594 ) );
  ADD32 \position1/sub_216_I2/U2_22  ( .A(\position1/N1568 ), .B(n269), .CI(
        \position1/sub_216_I2/carry [22]), .CO(
        \position1/sub_216_I2/carry [23]), .S(\position1/N1595 ) );
  ADD32 \position1/sub_216_I2/U2_23  ( .A(\position1/N1569 ), .B(n300), .CI(
        \position1/sub_216_I2/carry [23]), .CO(
        \position1/sub_216_I2/carry [24]), .S(\position1/N1596 ) );
  ADD32 \position1/sub_216_I3/U2_7  ( .A(n1298), .B(n36), .CI(
        \position1/sub_216_I3/carry [7]), .CO(\position1/sub_216_I3/carry [8]), 
        .S(\position1/N1632 ) );
  ADD32 \position1/sub_216_I3/U2_8  ( .A(n1296), .B(n245), .CI(
        \position1/sub_216_I3/carry [8]), .CO(\position1/sub_216_I3/carry [9]), 
        .S(\position1/N1633 ) );
  ADD32 \position1/sub_216_I3/U2_9  ( .A(n1293), .B(n246), .CI(
        \position1/sub_216_I3/carry [9]), .CO(\position1/sub_216_I3/carry [10]), .S(\position1/N1634 ) );
  ADD32 \position1/sub_216_I3/U2_10  ( .A(n1291), .B(n248), .CI(
        \position1/sub_216_I3/carry [10]), .CO(
        \position1/sub_216_I3/carry [11]), .S(\position1/N1635 ) );
  ADD32 \position1/sub_216_I3/U2_11  ( .A(n1288), .B(n47), .CI(
        \position1/sub_216_I3/carry [11]), .CO(
        \position1/sub_216_I3/carry [12]), .S(\position1/N1636 ) );
  ADD32 \position1/sub_216_I3/U2_12  ( .A(n1286), .B(n252), .CI(
        \position1/sub_216_I3/carry [12]), .CO(
        \position1/sub_216_I3/carry [13]), .S(\position1/N1637 ) );
  ADD32 \position1/sub_216_I3/U2_13  ( .A(n1284), .B(n254), .CI(
        \position1/sub_216_I3/carry [13]), .CO(
        \position1/sub_216_I3/carry [14]), .S(\position1/N1638 ) );
  ADD32 \position1/sub_216_I3/U2_14  ( .A(n1282), .B(n284), .CI(
        \position1/sub_216_I3/carry [14]), .CO(
        \position1/sub_216_I3/carry [15]), .S(\position1/N1639 ) );
  ADD32 \position1/sub_216_I3/U2_15  ( .A(n1280), .B(n286), .CI(
        \position1/sub_216_I3/carry [15]), .CO(
        \position1/sub_216_I3/carry [16]), .S(\position1/N1640 ) );
  ADD32 \position1/sub_216_I3/U2_16  ( .A(n1278), .B(n259), .CI(
        \position1/sub_216_I3/carry [16]), .CO(
        \position1/sub_216_I3/carry [17]), .S(\position1/N1641 ) );
  ADD32 \position1/sub_216_I3/U2_17  ( .A(n1276), .B(n261), .CI(
        \position1/sub_216_I3/carry [17]), .CO(
        \position1/sub_216_I3/carry [18]), .S(\position1/N1642 ) );
  ADD32 \position1/sub_216_I3/U2_18  ( .A(n1274), .B(n292), .CI(
        \position1/sub_216_I3/carry [18]), .CO(
        \position1/sub_216_I3/carry [19]), .S(\position1/N1643 ) );
  ADD32 \position1/sub_216_I3/U2_19  ( .A(n1272), .B(n265), .CI(
        \position1/sub_216_I3/carry [19]), .CO(
        \position1/sub_216_I3/carry [20]), .S(\position1/N1644 ) );
  ADD32 \position1/sub_216_I3/U2_20  ( .A(n1270), .B(n267), .CI(
        \position1/sub_216_I3/carry [20]), .CO(
        \position1/sub_216_I3/carry [21]), .S(\position1/N1645 ) );
  ADD32 \position1/sub_216_I3/U2_21  ( .A(n1268), .B(n67), .CI(
        \position1/sub_216_I3/carry [21]), .CO(
        \position1/sub_216_I3/carry [22]), .S(\position1/N1646 ) );
  ADD32 \position1/sub_216_I3/U2_22  ( .A(n1267), .B(n44), .CI(
        \position1/sub_216_I3/carry [22]), .CO(
        \position1/sub_216_I3/carry [23]), .S(\position1/N1647 ) );
  ADD32 \position1/sub_216_I3/U2_23  ( .A(n1266), .B(n587), .CI(
        \position1/sub_216_I3/carry [23]), .CO(
        \position1/sub_216_I3/carry [24]), .S(\position1/N1648 ) );
  ADD32 \position1/sub_216_I4/U2_6  ( .A(\position1/N1656 ), .B(n36), .CI(
        \position1/sub_216_I4/carry [6]), .CO(\position1/sub_216_I4/carry [7]), 
        .S(\position1/N1683 ) );
  ADD32 \position1/sub_216_I4/U2_7  ( .A(\position1/N1657 ), .B(n66), .CI(
        \position1/sub_216_I4/carry [7]), .CO(\position1/sub_216_I4/carry [8]), 
        .S(\position1/N1684 ) );
  ADD32 \position1/sub_216_I4/U2_8  ( .A(\position1/N1658 ), .B(n37), .CI(
        \position1/sub_216_I4/carry [8]), .CO(\position1/sub_216_I4/carry [9]), 
        .S(\position1/N1685 ) );
  ADD32 \position1/sub_216_I4/U2_9  ( .A(\position1/N1659 ), .B(n276), .CI(
        \position1/sub_216_I4/carry [9]), .CO(\position1/sub_216_I4/carry [10]), .S(\position1/N1686 ) );
  ADD32 \position1/sub_216_I4/U2_10  ( .A(\position1/N1660 ), .B(n250), .CI(
        \position1/sub_216_I4/carry [10]), .CO(
        \position1/sub_216_I4/carry [11]), .S(\position1/N1687 ) );
  ADD32 \position1/sub_216_I4/U2_11  ( .A(\position1/N1661 ), .B(n280), .CI(
        \position1/sub_216_I4/carry [11]), .CO(
        \position1/sub_216_I4/carry [12]), .S(\position1/N1688 ) );
  ADD32 \position1/sub_216_I4/U2_12  ( .A(\position1/N1662 ), .B(n100), .CI(
        \position1/sub_216_I4/carry [12]), .CO(
        \position1/sub_216_I4/carry [13]), .S(\position1/N1689 ) );
  ADD32 \position1/sub_216_I4/U2_13  ( .A(\position1/N1663 ), .B(n256), .CI(
        \position1/sub_216_I4/carry [13]), .CO(
        \position1/sub_216_I4/carry [14]), .S(\position1/N1690 ) );
  ADD32 \position1/sub_216_I4/U2_14  ( .A(\position1/N1664 ), .B(n35), .CI(
        \position1/sub_216_I4/carry [14]), .CO(
        \position1/sub_216_I4/carry [15]), .S(\position1/N1691 ) );
  ADD32 \position1/sub_216_I4/U2_15  ( .A(\position1/N1665 ), .B(n288), .CI(
        \position1/sub_216_I4/carry [15]), .CO(
        \position1/sub_216_I4/carry [16]), .S(\position1/N1692 ) );
  ADD32 \position1/sub_216_I4/U2_16  ( .A(\position1/N1666 ), .B(n38), .CI(
        \position1/sub_216_I4/carry [16]), .CO(
        \position1/sub_216_I4/carry [17]), .S(\position1/N1693 ) );
  ADD32 \position1/sub_216_I4/U2_17  ( .A(\position1/N1667 ), .B(n263), .CI(
        \position1/sub_216_I4/carry [17]), .CO(
        \position1/sub_216_I4/carry [18]), .S(\position1/N1694 ) );
  ADD32 \position1/sub_216_I4/U2_18  ( .A(\position1/N1668 ), .B(n39), .CI(
        \position1/sub_216_I4/carry [18]), .CO(
        \position1/sub_216_I4/carry [19]), .S(\position1/N1695 ) );
  ADD32 \position1/sub_216_I4/U2_19  ( .A(\position1/N1669 ), .B(n296), .CI(
        \position1/sub_216_I4/carry [19]), .CO(
        \position1/sub_216_I4/carry [20]), .S(\position1/N1696 ) );
  ADD32 \position1/sub_216_I4/U2_20  ( .A(\position1/N1670 ), .B(n298), .CI(
        \position1/sub_216_I4/carry [20]), .CO(
        \position1/sub_216_I4/carry [21]), .S(\position1/N1697 ) );
  ADD32 \position1/sub_216_I4/U2_21  ( .A(\position1/N1671 ), .B(n300), .CI(
        \position1/sub_216_I4/carry [21]), .CO(
        \position1/sub_216_I4/carry [22]), .S(\position1/N1698 ) );
  ADD32 \position1/sub_216_I4/U2_22  ( .A(\position1/N1672 ), .B(n587), .CI(
        \position1/sub_216_I4/carry [22]), .CO(
        \position1/sub_216_I4/carry [23]), .S(\position1/N1699 ) );
  ADD32 \position1/sub_216_I5/U2_5  ( .A(n1237), .B(n36), .CI(
        \position1/sub_216_I5/carry [5]), .CO(\position1/sub_216_I5/carry [6]), 
        .S(\position1/N1734 ) );
  ADD32 \position1/sub_216_I5/U2_6  ( .A(n1235), .B(n245), .CI(
        \position1/sub_216_I5/carry [6]), .CO(\position1/sub_216_I5/carry [7]), 
        .S(\position1/N1735 ) );
  ADD32 \position1/sub_216_I5/U2_7  ( .A(n1233), .B(n246), .CI(
        \position1/sub_216_I5/carry [7]), .CO(\position1/sub_216_I5/carry [8]), 
        .S(\position1/N1736 ) );
  ADD32 \position1/sub_216_I5/U2_8  ( .A(n1231), .B(n248), .CI(
        \position1/sub_216_I5/carry [8]), .CO(\position1/sub_216_I5/carry [9]), 
        .S(\position1/N1737 ) );
  ADD32 \position1/sub_216_I5/U2_9  ( .A(n1229), .B(n47), .CI(
        \position1/sub_216_I5/carry [9]), .CO(\position1/sub_216_I5/carry [10]), .S(\position1/N1738 ) );
  ADD32 \position1/sub_216_I5/U2_10  ( .A(n1228), .B(n252), .CI(
        \position1/sub_216_I5/carry [10]), .CO(
        \position1/sub_216_I5/carry [11]), .S(\position1/N1739 ) );
  ADD32 \position1/sub_216_I5/U2_11  ( .A(n1226), .B(n100), .CI(
        \position1/sub_216_I5/carry [11]), .CO(
        \position1/sub_216_I5/carry [12]), .S(\position1/N1740 ) );
  ADD32 \position1/sub_216_I5/U2_12  ( .A(n1225), .B(n284), .CI(
        \position1/sub_216_I5/carry [12]), .CO(
        \position1/sub_216_I5/carry [13]), .S(\position1/N1741 ) );
  ADD32 \position1/sub_216_I5/U2_13  ( .A(n1224), .B(n35), .CI(
        \position1/sub_216_I5/carry [13]), .CO(
        \position1/sub_216_I5/carry [14]), .S(\position1/N1742 ) );
  ADD32 \position1/sub_216_I5/U2_14  ( .A(n1223), .B(n259), .CI(
        \position1/sub_216_I5/carry [14]), .CO(
        \position1/sub_216_I5/carry [15]), .S(\position1/N1743 ) );
  ADD32 \position1/sub_216_I5/U2_15  ( .A(n1222), .B(n261), .CI(
        \position1/sub_216_I5/carry [15]), .CO(
        \position1/sub_216_I5/carry [16]), .S(\position1/N1744 ) );
  ADD32 \position1/sub_216_I5/U2_16  ( .A(n1221), .B(n292), .CI(
        \position1/sub_216_I5/carry [16]), .CO(
        \position1/sub_216_I5/carry [17]), .S(\position1/N1745 ) );
  ADD32 \position1/sub_216_I5/U2_17  ( .A(n1220), .B(n265), .CI(
        \position1/sub_216_I5/carry [17]), .CO(
        \position1/sub_216_I5/carry [18]), .S(\position1/N1746 ) );
  ADD32 \position1/sub_216_I5/U2_18  ( .A(n1219), .B(n267), .CI(
        \position1/sub_216_I5/carry [18]), .CO(
        \position1/sub_216_I5/carry [19]), .S(\position1/N1747 ) );
  ADD32 \position1/sub_216_I5/U2_19  ( .A(n1218), .B(n67), .CI(
        \position1/sub_216_I5/carry [19]), .CO(
        \position1/sub_216_I5/carry [20]), .S(\position1/N1748 ) );
  ADD32 \position1/sub_216_I5/U2_20  ( .A(n1217), .B(n44), .CI(
        \position1/sub_216_I5/carry [20]), .CO(
        \position1/sub_216_I5/carry [21]), .S(\position1/N1749 ) );
  ADD32 \position1/sub_216_I5/U2_21  ( .A(n1216), .B(n588), .CI(
        \position1/sub_216_I5/carry [21]), .CO(
        \position1/sub_216_I5/carry [22]), .S(\position1/N1750 ) );
  ADD32 \position1/sub_216_I6/U2_4  ( .A(n1207), .B(n36), .CI(
        \position1/sub_216_I6/carry [4]), .CO(\position1/sub_216_I6/carry [5]), 
        .S(\position1/N1785 ) );
  ADD32 \position1/sub_216_I6/U2_5  ( .A(n1206), .B(n66), .CI(
        \position1/sub_216_I6/carry [5]), .CO(\position1/sub_216_I6/carry [6]), 
        .S(\position1/N1786 ) );
  ADD32 \position1/sub_216_I6/U2_6  ( .A(n1205), .B(n37), .CI(
        \position1/sub_216_I6/carry [6]), .CO(\position1/sub_216_I6/carry [7]), 
        .S(\position1/N1787 ) );
  ADD32 \position1/sub_216_I6/U2_7  ( .A(n1204), .B(n276), .CI(
        \position1/sub_216_I6/carry [7]), .CO(\position1/sub_216_I6/carry [8]), 
        .S(\position1/N1788 ) );
  ADD32 \position1/sub_216_I6/U2_8  ( .A(n1203), .B(n47), .CI(
        \position1/sub_216_I6/carry [8]), .CO(\position1/sub_216_I6/carry [9]), 
        .S(\position1/N1789 ) );
  ADD32 \position1/sub_216_I6/U2_9  ( .A(n1202), .B(n280), .CI(
        \position1/sub_216_I6/carry [9]), .CO(\position1/sub_216_I6/carry [10]), .S(\position1/N1790 ) );
  ADD32 \position1/sub_216_I6/U2_10  ( .A(n1201), .B(n100), .CI(
        \position1/sub_216_I6/carry [10]), .CO(
        \position1/sub_216_I6/carry [11]), .S(\position1/N1791 ) );
  ADD32 \position1/sub_216_I6/U2_11  ( .A(n1200), .B(n256), .CI(
        \position1/sub_216_I6/carry [11]), .CO(
        \position1/sub_216_I6/carry [12]), .S(\position1/N1792 ) );
  ADD32 \position1/sub_216_I6/U2_12  ( .A(n1199), .B(n35), .CI(
        \position1/sub_216_I6/carry [12]), .CO(
        \position1/sub_216_I6/carry [13]), .S(\position1/N1793 ) );
  ADD32 \position1/sub_216_I6/U2_13  ( .A(n1198), .B(n288), .CI(
        \position1/sub_216_I6/carry [13]), .CO(
        \position1/sub_216_I6/carry [14]), .S(\position1/N1794 ) );
  ADD32 \position1/sub_216_I6/U2_14  ( .A(n1197), .B(n38), .CI(
        \position1/sub_216_I6/carry [14]), .CO(
        \position1/sub_216_I6/carry [15]), .S(\position1/N1795 ) );
  ADD32 \position1/sub_216_I6/U2_15  ( .A(n1196), .B(n263), .CI(
        \position1/sub_216_I6/carry [15]), .CO(
        \position1/sub_216_I6/carry [16]), .S(\position1/N1796 ) );
  ADD32 \position1/sub_216_I6/U2_16  ( .A(n1195), .B(n39), .CI(
        \position1/sub_216_I6/carry [16]), .CO(
        \position1/sub_216_I6/carry [17]), .S(\position1/N1797 ) );
  ADD32 \position1/sub_216_I6/U2_17  ( .A(n1194), .B(n296), .CI(
        \position1/sub_216_I6/carry [17]), .CO(
        \position1/sub_216_I6/carry [18]), .S(\position1/N1798 ) );
  ADD32 \position1/sub_216_I6/U2_18  ( .A(n1192), .B(n67), .CI(
        \position1/sub_216_I6/carry [18]), .CO(
        \position1/sub_216_I6/carry [19]), .S(\position1/N1799 ) );
  ADD32 \position1/sub_216_I6/U2_19  ( .A(n1191), .B(n300), .CI(
        \position1/sub_216_I6/carry [19]), .CO(
        \position1/sub_216_I6/carry [20]), .S(\position1/N1800 ) );
  ADD32 \position1/sub_216_I6/U2_20  ( .A(n1189), .B(n588), .CI(
        \position1/sub_216_I6/carry [20]), .CO(
        \position1/sub_216_I6/carry [21]), .S(\position1/N1801 ) );
  ADD32 \position1/sub_216_I7/U2_3  ( .A(n1180), .B(n628), .CI(
        \position1/sub_216_I7/carry [3]), .CO(\position1/sub_216_I7/carry [4]), 
        .S(\position1/N1836 ) );
  ADD32 \position1/sub_216_I7/U2_4  ( .A(n1179), .B(n66), .CI(
        \position1/sub_216_I7/carry [4]), .CO(\position1/sub_216_I7/carry [5]), 
        .S(\position1/N1837 ) );
  ADD32 \position1/sub_216_I7/U2_5  ( .A(n1178), .B(n37), .CI(
        \position1/sub_216_I7/carry [5]), .CO(\position1/sub_216_I7/carry [6]), 
        .S(\position1/N1838 ) );
  ADD32 \position1/sub_216_I7/U2_6  ( .A(n1177), .B(n248), .CI(
        \position1/sub_216_I7/carry [6]), .CO(\position1/sub_216_I7/carry [7]), 
        .S(\position1/N1839 ) );
  ADD32 \position1/sub_216_I7/U2_7  ( .A(n1176), .B(n47), .CI(
        \position1/sub_216_I7/carry [7]), .CO(\position1/sub_216_I7/carry [8]), 
        .S(\position1/N1840 ) );
  ADD32 \position1/sub_216_I7/U2_8  ( .A(n1175), .B(n252), .CI(
        \position1/sub_216_I7/carry [8]), .CO(\position1/sub_216_I7/carry [9]), 
        .S(\position1/N1841 ) );
  ADD32 \position1/sub_216_I7/U2_9  ( .A(n1174), .B(n100), .CI(
        \position1/sub_216_I7/carry [9]), .CO(\position1/sub_216_I7/carry [10]), .S(\position1/N1842 ) );
  ADD32 \position1/sub_216_I7/U2_10  ( .A(n1173), .B(n284), .CI(
        \position1/sub_216_I7/carry [10]), .CO(
        \position1/sub_216_I7/carry [11]), .S(\position1/N1843 ) );
  ADD32 \position1/sub_216_I7/U2_11  ( .A(n1172), .B(n35), .CI(
        \position1/sub_216_I7/carry [11]), .CO(
        \position1/sub_216_I7/carry [12]), .S(\position1/N1844 ) );
  ADD32 \position1/sub_216_I7/U2_12  ( .A(n1171), .B(n259), .CI(
        \position1/sub_216_I7/carry [12]), .CO(
        \position1/sub_216_I7/carry [13]), .S(\position1/N1845 ) );
  ADD32 \position1/sub_216_I7/U2_13  ( .A(n1170), .B(n38), .CI(
        \position1/sub_216_I7/carry [13]), .CO(
        \position1/sub_216_I7/carry [14]), .S(\position1/N1846 ) );
  ADD32 \position1/sub_216_I7/U2_14  ( .A(n1169), .B(n292), .CI(
        \position1/sub_216_I7/carry [14]), .CO(
        \position1/sub_216_I7/carry [15]), .S(\position1/N1847 ) );
  ADD32 \position1/sub_216_I7/U2_15  ( .A(n1168), .B(n39), .CI(
        \position1/sub_216_I7/carry [15]), .CO(
        \position1/sub_216_I7/carry [16]), .S(\position1/N1848 ) );
  ADD32 \position1/sub_216_I7/U2_16  ( .A(n1167), .B(n296), .CI(
        \position1/sub_216_I7/carry [16]), .CO(
        \position1/sub_216_I7/carry [17]), .S(\position1/N1849 ) );
  ADD32 \position1/sub_216_I7/U2_17  ( .A(n1166), .B(n67), .CI(
        \position1/sub_216_I7/carry [17]), .CO(
        \position1/sub_216_I7/carry [18]), .S(\position1/N1850 ) );
  ADD32 \position1/sub_216_I7/U2_18  ( .A(n1165), .B(n44), .CI(
        \position1/sub_216_I7/carry [18]), .CO(
        \position1/sub_216_I7/carry [19]), .S(\position1/N1851 ) );
  ADD32 \position1/sub_216_I7/U2_19  ( .A(n1164), .B(n588), .CI(
        \position1/sub_216_I7/carry [19]), .CO(
        \position1/sub_216_I7/carry [20]), .S(\position1/N1852 ) );
  ADD32 \position1/sub_216_I8/U2_2  ( .A(n1155), .B(n36), .CI(
        \position1/sub_216_I8/carry [2]), .CO(\position1/sub_216_I8/carry [3]), 
        .S(\position1/N1887 ) );
  ADD32 \position1/sub_216_I8/U2_3  ( .A(n1153), .B(n66), .CI(
        \position1/sub_216_I8/carry [3]), .CO(\position1/sub_216_I8/carry [4]), 
        .S(\position1/N1888 ) );
  ADD32 \position1/sub_216_I8/U2_4  ( .A(n1152), .B(n37), .CI(
        \position1/sub_216_I8/carry [4]), .CO(\position1/sub_216_I8/carry [5]), 
        .S(\position1/N1889 ) );
  ADD32 \position1/sub_216_I8/U2_5  ( .A(n1150), .B(n276), .CI(
        \position1/sub_216_I8/carry [5]), .CO(\position1/sub_216_I8/carry [6]), 
        .S(\position1/N1890 ) );
  ADD32 \position1/sub_216_I8/U2_6  ( .A(n1149), .B(n47), .CI(
        \position1/sub_216_I8/carry [6]), .CO(\position1/sub_216_I8/carry [7]), 
        .S(\position1/N1891 ) );
  ADD32 \position1/sub_216_I8/U2_7  ( .A(n1147), .B(n280), .CI(
        \position1/sub_216_I8/carry [7]), .CO(\position1/sub_216_I8/carry [8]), 
        .S(\position1/N1892 ) );
  ADD32 \position1/sub_216_I8/U2_8  ( .A(n1146), .B(n100), .CI(
        \position1/sub_216_I8/carry [8]), .CO(\position1/sub_216_I8/carry [9]), 
        .S(\position1/N1893 ) );
  ADD32 \position1/sub_216_I8/U2_9  ( .A(n1144), .B(n284), .CI(
        \position1/sub_216_I8/carry [9]), .CO(\position1/sub_216_I8/carry [10]), .S(\position1/N1894 ) );
  ADD32 \position1/sub_216_I8/U2_10  ( .A(n1143), .B(n35), .CI(
        \position1/sub_216_I8/carry [10]), .CO(
        \position1/sub_216_I8/carry [11]), .S(\position1/N1895 ) );
  ADD32 \position1/sub_216_I8/U2_11  ( .A(n1142), .B(n288), .CI(
        \position1/sub_216_I8/carry [11]), .CO(
        \position1/sub_216_I8/carry [12]), .S(\position1/N1896 ) );
  ADD32 \position1/sub_216_I8/U2_12  ( .A(n1140), .B(n38), .CI(
        \position1/sub_216_I8/carry [12]), .CO(
        \position1/sub_216_I8/carry [13]), .S(\position1/N1897 ) );
  ADD32 \position1/sub_216_I8/U2_13  ( .A(n1138), .B(n292), .CI(
        \position1/sub_216_I8/carry [13]), .CO(
        \position1/sub_216_I8/carry [14]), .S(\position1/N1898 ) );
  ADD32 \position1/sub_216_I8/U2_14  ( .A(n1137), .B(n39), .CI(
        \position1/sub_216_I8/carry [14]), .CO(
        \position1/sub_216_I8/carry [15]), .S(\position1/N1899 ) );
  ADD32 \position1/sub_216_I8/U2_15  ( .A(n1135), .B(n296), .CI(
        \position1/sub_216_I8/carry [15]), .CO(
        \position1/sub_216_I8/carry [16]), .S(\position1/N1900 ) );
  ADD32 \position1/sub_216_I8/U2_16  ( .A(n1134), .B(n67), .CI(
        \position1/sub_216_I8/carry [16]), .CO(
        \position1/sub_216_I8/carry [17]), .S(\position1/N1901 ) );
  ADD32 \position1/sub_216_I8/U2_17  ( .A(n1133), .B(n44), .CI(
        \position1/sub_216_I8/carry [17]), .CO(
        \position1/sub_216_I8/carry [18]), .S(\position1/N1902 ) );
  ADD32 \position1/sub_216_I8/U2_18  ( .A(n1132), .B(n588), .CI(
        \position1/sub_216_I8/carry [18]), .CO(
        \position1/sub_216_I8/carry [19]), .S(\position1/N1903 ) );
  ADD32 \position1/sub_226/U2_9  ( .A(\position1/y_sum [9]), .B(n36), .CI(
        \position1/sub_226/carry [9]), .CO(\position1/sub_226/carry [10]), .S(
        \position1/N1947 ) );
  ADD32 \position1/sub_226/U2_10  ( .A(\position1/y_sum [10]), .B(n66), .CI(
        \position1/sub_226/carry [10]), .CO(\position1/sub_226/carry [11]), 
        .S(\position1/N1948 ) );
  ADD32 \position1/sub_226/U2_11  ( .A(\position1/y_sum [11]), .B(n37), .CI(
        \position1/sub_226/carry [11]), .CO(\position1/sub_226/carry [12]), 
        .S(\position1/N1949 ) );
  ADD32 \position1/sub_226/U2_12  ( .A(\position1/y_sum [12]), .B(n41), .CI(
        \position1/sub_226/carry [12]), .CO(\position1/sub_226/carry [13]), 
        .S(\position1/N1950 ) );
  ADD32 \position1/sub_226/U2_13  ( .A(\position1/y_sum [13]), .B(n47), .CI(
        \position1/sub_226/carry [13]), .CO(\position1/sub_226/carry [14]), 
        .S(\position1/N1951 ) );
  ADD32 \position1/sub_226/U2_14  ( .A(\position1/y_sum [14]), .B(n45), .CI(
        \position1/sub_226/carry [14]), .CO(\position1/sub_226/carry [15]), 
        .S(\position1/N1952 ) );
  ADD32 \position1/sub_226/U2_15  ( .A(\position1/y_sum [15]), .B(n100), .CI(
        \position1/sub_226/carry [15]), .CO(\position1/sub_226/carry [16]), 
        .S(\position1/N1953 ) );
  ADD32 \position1/sub_226/U2_16  ( .A(\position1/y_sum [16]), .B(n40), .CI(
        \position1/sub_226/carry [16]), .CO(\position1/sub_226/carry [17]), 
        .S(\position1/N1954 ) );
  ADD32 \position1/sub_226/U2_17  ( .A(\position1/y_sum [17]), .B(n35), .CI(
        \position1/sub_226/carry [17]), .CO(\position1/sub_226/carry [18]), 
        .S(\position1/N1955 ) );
  ADD32 \position1/sub_226/U2_18  ( .A(\position1/y_sum [18]), .B(n288), .CI(
        \position1/sub_226/carry [18]), .CO(\position1/sub_226/carry [19]), 
        .S(\position1/N1956 ) );
  ADD32 \position1/sub_226/U2_19  ( .A(\position1/y_sum [19]), .B(n38), .CI(
        \position1/sub_226/carry [19]), .CO(\position1/sub_226/carry [20]), 
        .S(\position1/N1957 ) );
  ADD32 \position1/sub_226/U2_20  ( .A(\position1/y_sum [20]), .B(n43), .CI(
        \position1/sub_226/carry [20]), .CO(\position1/sub_226/carry [21]), 
        .S(\position1/N1958 ) );
  ADD32 \position1/sub_226/U2_21  ( .A(\position1/y_sum [21]), .B(n39), .CI(
        \position1/sub_226/carry [21]), .CO(\position1/sub_226/carry [22]), 
        .S(\position1/N1959 ) );
  ADD32 \position1/sub_226/U2_22  ( .A(\position1/y_sum [22]), .B(n42), .CI(
        \position1/sub_226/carry [22]), .CO(\position1/sub_226/carry [23]), 
        .S(\position1/N1960 ) );
  ADD32 \position1/sub_226/U2_23  ( .A(\position1/y_sum [23]), .B(n67), .CI(
        \position1/sub_226/carry [23]), .CO(\position1/sub_226/carry [24]), 
        .S(\position1/N1961 ) );
  ADD32 \position1/sub_226_I2/U2_8  ( .A(\position1/N1971 ), .B(n628), .CI(
        \position1/sub_226_I2/carry [8]), .CO(\position1/sub_226_I2/carry [9]), 
        .S(\position1/N1998 ) );
  ADD32 \position1/sub_226_I2/U2_9  ( .A(\position1/N1972 ), .B(n66), .CI(
        \position1/sub_226_I2/carry [9]), .CO(\position1/sub_226_I2/carry [10]), .S(\position1/N1999 ) );
  ADD32 \position1/sub_226_I2/U2_10  ( .A(\position1/N1973 ), .B(n37), .CI(
        \position1/sub_226_I2/carry [10]), .CO(
        \position1/sub_226_I2/carry [11]), .S(\position1/N2000 ) );
  ADD32 \position1/sub_226_I2/U2_11  ( .A(\position1/N1974 ), .B(n41), .CI(
        \position1/sub_226_I2/carry [11]), .CO(
        \position1/sub_226_I2/carry [12]), .S(\position1/N2001 ) );
  ADD32 \position1/sub_226_I2/U2_12  ( .A(\position1/N1975 ), .B(n47), .CI(
        \position1/sub_226_I2/carry [12]), .CO(
        \position1/sub_226_I2/carry [13]), .S(\position1/N2002 ) );
  ADD32 \position1/sub_226_I2/U2_13  ( .A(\position1/N1976 ), .B(n45), .CI(
        \position1/sub_226_I2/carry [13]), .CO(
        \position1/sub_226_I2/carry [14]), .S(\position1/N2003 ) );
  ADD32 \position1/sub_226_I2/U2_14  ( .A(\position1/N1977 ), .B(n100), .CI(
        \position1/sub_226_I2/carry [14]), .CO(
        \position1/sub_226_I2/carry [15]), .S(\position1/N2004 ) );
  ADD32 \position1/sub_226_I2/U2_15  ( .A(\position1/N1978 ), .B(n40), .CI(
        \position1/sub_226_I2/carry [15]), .CO(
        \position1/sub_226_I2/carry [16]), .S(\position1/N2005 ) );
  ADD32 \position1/sub_226_I2/U2_16  ( .A(\position1/N1979 ), .B(n35), .CI(
        \position1/sub_226_I2/carry [16]), .CO(
        \position1/sub_226_I2/carry [17]), .S(\position1/N2006 ) );
  ADD32 \position1/sub_226_I2/U2_17  ( .A(\position1/N1980 ), .B(n46), .CI(
        \position1/sub_226_I2/carry [17]), .CO(
        \position1/sub_226_I2/carry [18]), .S(\position1/N2007 ) );
  ADD32 \position1/sub_226_I2/U2_18  ( .A(\position1/N1981 ), .B(n38), .CI(
        \position1/sub_226_I2/carry [18]), .CO(
        \position1/sub_226_I2/carry [19]), .S(\position1/N2008 ) );
  ADD32 \position1/sub_226_I2/U2_19  ( .A(\position1/N1982 ), .B(n43), .CI(
        \position1/sub_226_I2/carry [19]), .CO(
        \position1/sub_226_I2/carry [20]), .S(\position1/N2009 ) );
  ADD32 \position1/sub_226_I2/U2_20  ( .A(\position1/N1983 ), .B(n39), .CI(
        \position1/sub_226_I2/carry [20]), .CO(
        \position1/sub_226_I2/carry [21]), .S(\position1/N2010 ) );
  ADD32 \position1/sub_226_I2/U2_21  ( .A(\position1/N1984 ), .B(n42), .CI(
        \position1/sub_226_I2/carry [21]), .CO(
        \position1/sub_226_I2/carry [22]), .S(\position1/N2011 ) );
  ADD32 \position1/sub_226_I2/U2_22  ( .A(\position1/N1985 ), .B(n67), .CI(
        \position1/sub_226_I2/carry [22]), .CO(
        \position1/sub_226_I2/carry [23]), .S(\position1/N2012 ) );
  ADD32 \position1/sub_226_I2/U2_23  ( .A(\position1/N1986 ), .B(n44), .CI(
        \position1/sub_226_I2/carry [23]), .CO(
        \position1/sub_226_I2/carry [24]), .S(\position1/N2013 ) );
  ADD32 \position1/sub_226_I3/U2_7  ( .A(n1079), .B(n36), .CI(
        \position1/sub_226_I3/carry [7]), .CO(\position1/sub_226_I3/carry [8]), 
        .S(\position1/N2049 ) );
  ADD32 \position1/sub_226_I3/U2_8  ( .A(n1077), .B(n66), .CI(
        \position1/sub_226_I3/carry [8]), .CO(\position1/sub_226_I3/carry [9]), 
        .S(\position1/N2050 ) );
  ADD32 \position1/sub_226_I3/U2_9  ( .A(n1074), .B(n37), .CI(
        \position1/sub_226_I3/carry [9]), .CO(\position1/sub_226_I3/carry [10]), .S(\position1/N2051 ) );
  ADD32 \position1/sub_226_I3/U2_10  ( .A(n1072), .B(n41), .CI(
        \position1/sub_226_I3/carry [10]), .CO(
        \position1/sub_226_I3/carry [11]), .S(\position1/N2052 ) );
  ADD32 \position1/sub_226_I3/U2_11  ( .A(n1069), .B(n47), .CI(
        \position1/sub_226_I3/carry [11]), .CO(
        \position1/sub_226_I3/carry [12]), .S(\position1/N2053 ) );
  ADD32 \position1/sub_226_I3/U2_12  ( .A(n1067), .B(n45), .CI(
        \position1/sub_226_I3/carry [12]), .CO(
        \position1/sub_226_I3/carry [13]), .S(\position1/N2054 ) );
  ADD32 \position1/sub_226_I3/U2_13  ( .A(n1065), .B(n100), .CI(
        \position1/sub_226_I3/carry [13]), .CO(
        \position1/sub_226_I3/carry [14]), .S(\position1/N2055 ) );
  ADD32 \position1/sub_226_I3/U2_14  ( .A(n1063), .B(n40), .CI(
        \position1/sub_226_I3/carry [14]), .CO(
        \position1/sub_226_I3/carry [15]), .S(\position1/N2056 ) );
  ADD32 \position1/sub_226_I3/U2_15  ( .A(n1061), .B(n35), .CI(
        \position1/sub_226_I3/carry [15]), .CO(
        \position1/sub_226_I3/carry [16]), .S(\position1/N2057 ) );
  ADD32 \position1/sub_226_I3/U2_16  ( .A(n1059), .B(n46), .CI(
        \position1/sub_226_I3/carry [16]), .CO(
        \position1/sub_226_I3/carry [17]), .S(\position1/N2058 ) );
  ADD32 \position1/sub_226_I3/U2_17  ( .A(n1057), .B(n38), .CI(
        \position1/sub_226_I3/carry [17]), .CO(
        \position1/sub_226_I3/carry [18]), .S(\position1/N2059 ) );
  ADD32 \position1/sub_226_I3/U2_18  ( .A(n1055), .B(n43), .CI(
        \position1/sub_226_I3/carry [18]), .CO(
        \position1/sub_226_I3/carry [19]), .S(\position1/N2060 ) );
  ADD32 \position1/sub_226_I3/U2_19  ( .A(n1053), .B(n39), .CI(
        \position1/sub_226_I3/carry [19]), .CO(
        \position1/sub_226_I3/carry [20]), .S(\position1/N2061 ) );
  ADD32 \position1/sub_226_I3/U2_20  ( .A(n1051), .B(n42), .CI(
        \position1/sub_226_I3/carry [20]), .CO(
        \position1/sub_226_I3/carry [21]), .S(\position1/N2062 ) );
  ADD32 \position1/sub_226_I3/U2_21  ( .A(n1049), .B(n67), .CI(
        \position1/sub_226_I3/carry [21]), .CO(
        \position1/sub_226_I3/carry [22]), .S(\position1/N2063 ) );
  ADD32 \position1/sub_226_I3/U2_22  ( .A(n1048), .B(n44), .CI(
        \position1/sub_226_I3/carry [22]), .CO(
        \position1/sub_226_I3/carry [23]), .S(\position1/N2064 ) );
  ADD32 \position1/sub_226_I3/U2_23  ( .A(n1047), .B(n589), .CI(
        \position1/sub_226_I3/carry [23]), .CO(
        \position1/sub_226_I3/carry [24]), .S(\position1/N2065 ) );
  ADD32 \position1/sub_226_I4/U2_6  ( .A(\position1/N2073 ), .B(n628), .CI(
        \position1/sub_226_I4/carry [6]), .CO(\position1/sub_226_I4/carry [7]), 
        .S(\position1/N2100 ) );
  ADD32 \position1/sub_226_I4/U2_7  ( .A(\position1/N2074 ), .B(n66), .CI(
        \position1/sub_226_I4/carry [7]), .CO(\position1/sub_226_I4/carry [8]), 
        .S(\position1/N2101 ) );
  ADD32 \position1/sub_226_I4/U2_8  ( .A(\position1/N2075 ), .B(n37), .CI(
        \position1/sub_226_I4/carry [8]), .CO(\position1/sub_226_I4/carry [9]), 
        .S(\position1/N2102 ) );
  ADD32 \position1/sub_226_I4/U2_9  ( .A(\position1/N2076 ), .B(n41), .CI(
        \position1/sub_226_I4/carry [9]), .CO(\position1/sub_226_I4/carry [10]), .S(\position1/N2103 ) );
  ADD32 \position1/sub_226_I4/U2_10  ( .A(\position1/N2077 ), .B(n47), .CI(
        \position1/sub_226_I4/carry [10]), .CO(
        \position1/sub_226_I4/carry [11]), .S(\position1/N2104 ) );
  ADD32 \position1/sub_226_I4/U2_11  ( .A(\position1/N2078 ), .B(n45), .CI(
        \position1/sub_226_I4/carry [11]), .CO(
        \position1/sub_226_I4/carry [12]), .S(\position1/N2105 ) );
  ADD32 \position1/sub_226_I4/U2_12  ( .A(\position1/N2079 ), .B(n100), .CI(
        \position1/sub_226_I4/carry [12]), .CO(
        \position1/sub_226_I4/carry [13]), .S(\position1/N2106 ) );
  ADD32 \position1/sub_226_I4/U2_13  ( .A(\position1/N2080 ), .B(n40), .CI(
        \position1/sub_226_I4/carry [13]), .CO(
        \position1/sub_226_I4/carry [14]), .S(\position1/N2107 ) );
  ADD32 \position1/sub_226_I4/U2_14  ( .A(\position1/N2081 ), .B(n35), .CI(
        \position1/sub_226_I4/carry [14]), .CO(
        \position1/sub_226_I4/carry [15]), .S(\position1/N2108 ) );
  ADD32 \position1/sub_226_I4/U2_15  ( .A(\position1/N2082 ), .B(n46), .CI(
        \position1/sub_226_I4/carry [15]), .CO(
        \position1/sub_226_I4/carry [16]), .S(\position1/N2109 ) );
  ADD32 \position1/sub_226_I4/U2_16  ( .A(\position1/N2083 ), .B(n38), .CI(
        \position1/sub_226_I4/carry [16]), .CO(
        \position1/sub_226_I4/carry [17]), .S(\position1/N2110 ) );
  ADD32 \position1/sub_226_I4/U2_17  ( .A(\position1/N2084 ), .B(n43), .CI(
        \position1/sub_226_I4/carry [17]), .CO(
        \position1/sub_226_I4/carry [18]), .S(\position1/N2111 ) );
  ADD32 \position1/sub_226_I4/U2_18  ( .A(\position1/N2085 ), .B(n39), .CI(
        \position1/sub_226_I4/carry [18]), .CO(
        \position1/sub_226_I4/carry [19]), .S(\position1/N2112 ) );
  ADD32 \position1/sub_226_I4/U2_19  ( .A(\position1/N2086 ), .B(n42), .CI(
        \position1/sub_226_I4/carry [19]), .CO(
        \position1/sub_226_I4/carry [20]), .S(\position1/N2113 ) );
  ADD32 \position1/sub_226_I4/U2_20  ( .A(\position1/N2087 ), .B(n67), .CI(
        \position1/sub_226_I4/carry [20]), .CO(
        \position1/sub_226_I4/carry [21]), .S(\position1/N2114 ) );
  ADD32 \position1/sub_226_I4/U2_21  ( .A(\position1/N2088 ), .B(n44), .CI(
        \position1/sub_226_I4/carry [21]), .CO(
        \position1/sub_226_I4/carry [22]), .S(\position1/N2115 ) );
  ADD32 \position1/sub_226_I4/U2_22  ( .A(\position1/N2089 ), .B(n589), .CI(
        \position1/sub_226_I4/carry [22]), .CO(
        \position1/sub_226_I4/carry [23]), .S(\position1/N2116 ) );
  ADD32 \position1/sub_226_I5/U2_5  ( .A(n1018), .B(n36), .CI(
        \position1/sub_226_I5/carry [5]), .CO(\position1/sub_226_I5/carry [6]), 
        .S(\position1/N2151 ) );
  ADD32 \position1/sub_226_I5/U2_6  ( .A(n1016), .B(n245), .CI(
        \position1/sub_226_I5/carry [6]), .CO(\position1/sub_226_I5/carry [7]), 
        .S(\position1/N2152 ) );
  ADD32 \position1/sub_226_I5/U2_7  ( .A(n1014), .B(n274), .CI(
        \position1/sub_226_I5/carry [7]), .CO(\position1/sub_226_I5/carry [8]), 
        .S(\position1/N2153 ) );
  ADD32 \position1/sub_226_I5/U2_8  ( .A(n1012), .B(n41), .CI(
        \position1/sub_226_I5/carry [8]), .CO(\position1/sub_226_I5/carry [9]), 
        .S(\position1/N2154 ) );
  ADD32 \position1/sub_226_I5/U2_9  ( .A(n1010), .B(n278), .CI(
        \position1/sub_226_I5/carry [9]), .CO(\position1/sub_226_I5/carry [10]), .S(\position1/N2155 ) );
  ADD32 \position1/sub_226_I5/U2_10  ( .A(n1009), .B(n45), .CI(
        \position1/sub_226_I5/carry [10]), .CO(
        \position1/sub_226_I5/carry [11]), .S(\position1/N2156 ) );
  ADD32 \position1/sub_226_I5/U2_11  ( .A(n1007), .B(n100), .CI(
        \position1/sub_226_I5/carry [11]), .CO(
        \position1/sub_226_I5/carry [12]), .S(\position1/N2157 ) );
  ADD32 \position1/sub_226_I5/U2_12  ( .A(n1006), .B(n40), .CI(
        \position1/sub_226_I5/carry [12]), .CO(
        \position1/sub_226_I5/carry [13]), .S(\position1/N2158 ) );
  ADD32 \position1/sub_226_I5/U2_13  ( .A(n1005), .B(n35), .CI(
        \position1/sub_226_I5/carry [13]), .CO(
        \position1/sub_226_I5/carry [14]), .S(\position1/N2159 ) );
  ADD32 \position1/sub_226_I5/U2_14  ( .A(n1004), .B(n46), .CI(
        \position1/sub_226_I5/carry [14]), .CO(
        \position1/sub_226_I5/carry [15]), .S(\position1/N2160 ) );
  ADD32 \position1/sub_226_I5/U2_15  ( .A(n1003), .B(n261), .CI(
        \position1/sub_226_I5/carry [15]), .CO(
        \position1/sub_226_I5/carry [16]), .S(\position1/N2161 ) );
  ADD32 \position1/sub_226_I5/U2_16  ( .A(n1002), .B(n292), .CI(
        \position1/sub_226_I5/carry [16]), .CO(
        \position1/sub_226_I5/carry [17]), .S(\position1/N2162 ) );
  ADD32 \position1/sub_226_I5/U2_17  ( .A(n1001), .B(n265), .CI(
        \position1/sub_226_I5/carry [17]), .CO(
        \position1/sub_226_I5/carry [18]), .S(\position1/N2163 ) );
  ADD32 \position1/sub_226_I5/U2_18  ( .A(n1000), .B(n267), .CI(
        \position1/sub_226_I5/carry [18]), .CO(
        \position1/sub_226_I5/carry [19]), .S(\position1/N2164 ) );
  ADD32 \position1/sub_226_I5/U2_19  ( .A(n999), .B(n269), .CI(
        \position1/sub_226_I5/carry [19]), .CO(
        \position1/sub_226_I5/carry [20]), .S(\position1/N2165 ) );
  ADD32 \position1/sub_226_I5/U2_20  ( .A(n998), .B(n300), .CI(
        \position1/sub_226_I5/carry [20]), .CO(
        \position1/sub_226_I5/carry [21]), .S(\position1/N2166 ) );
  ADD32 \position1/sub_226_I5/U2_21  ( .A(n997), .B(n589), .CI(
        \position1/sub_226_I5/carry [21]), .CO(
        \position1/sub_226_I5/carry [22]), .S(\position1/N2167 ) );
  ADD32 \position1/sub_226_I6/U2_4  ( .A(n988), .B(n36), .CI(
        \position1/sub_226_I6/carry [4]), .CO(\position1/sub_226_I6/carry [5]), 
        .S(\position1/N2202 ) );
  ADD32 \position1/sub_226_I6/U2_5  ( .A(n987), .B(n272), .CI(
        \position1/sub_226_I6/carry [5]), .CO(\position1/sub_226_I6/carry [6]), 
        .S(\position1/N2203 ) );
  ADD32 \position1/sub_226_I6/U2_6  ( .A(n986), .B(n246), .CI(
        \position1/sub_226_I6/carry [6]), .CO(\position1/sub_226_I6/carry [7]), 
        .S(\position1/N2204 ) );
  ADD32 \position1/sub_226_I6/U2_7  ( .A(n985), .B(n41), .CI(
        \position1/sub_226_I6/carry [7]), .CO(\position1/sub_226_I6/carry [8]), 
        .S(\position1/N2205 ) );
  ADD32 \position1/sub_226_I6/U2_8  ( .A(n984), .B(n250), .CI(
        \position1/sub_226_I6/carry [8]), .CO(\position1/sub_226_I6/carry [9]), 
        .S(\position1/N2206 ) );
  ADD32 \position1/sub_226_I6/U2_9  ( .A(n983), .B(n45), .CI(
        \position1/sub_226_I6/carry [9]), .CO(\position1/sub_226_I6/carry [10]), .S(\position1/N2207 ) );
  ADD32 \position1/sub_226_I6/U2_10  ( .A(n982), .B(n254), .CI(
        \position1/sub_226_I6/carry [10]), .CO(
        \position1/sub_226_I6/carry [11]), .S(\position1/N2208 ) );
  ADD32 \position1/sub_226_I6/U2_11  ( .A(n981), .B(n40), .CI(
        \position1/sub_226_I6/carry [11]), .CO(
        \position1/sub_226_I6/carry [12]), .S(\position1/N2209 ) );
  ADD32 \position1/sub_226_I6/U2_12  ( .A(n980), .B(n286), .CI(
        \position1/sub_226_I6/carry [12]), .CO(
        \position1/sub_226_I6/carry [13]), .S(\position1/N2210 ) );
  ADD32 \position1/sub_226_I6/U2_13  ( .A(n979), .B(n46), .CI(
        \position1/sub_226_I6/carry [13]), .CO(
        \position1/sub_226_I6/carry [14]), .S(\position1/N2211 ) );
  ADD32 \position1/sub_226_I6/U2_14  ( .A(n978), .B(n290), .CI(
        \position1/sub_226_I6/carry [14]), .CO(
        \position1/sub_226_I6/carry [15]), .S(\position1/N2212 ) );
  ADD32 \position1/sub_226_I6/U2_15  ( .A(n977), .B(n43), .CI(
        \position1/sub_226_I6/carry [15]), .CO(
        \position1/sub_226_I6/carry [16]), .S(\position1/N2213 ) );
  ADD32 \position1/sub_226_I6/U2_16  ( .A(n976), .B(n294), .CI(
        \position1/sub_226_I6/carry [16]), .CO(
        \position1/sub_226_I6/carry [17]), .S(\position1/N2214 ) );
  ADD32 \position1/sub_226_I6/U2_17  ( .A(n975), .B(n42), .CI(
        \position1/sub_226_I6/carry [17]), .CO(
        \position1/sub_226_I6/carry [18]), .S(\position1/N2215 ) );
  ADD32 \position1/sub_226_I6/U2_18  ( .A(n973), .B(n298), .CI(
        \position1/sub_226_I6/carry [18]), .CO(
        \position1/sub_226_I6/carry [19]), .S(\position1/N2216 ) );
  ADD32 \position1/sub_226_I6/U2_19  ( .A(n972), .B(n300), .CI(
        \position1/sub_226_I6/carry [19]), .CO(
        \position1/sub_226_I6/carry [20]), .S(\position1/N2217 ) );
  ADD32 \position1/sub_226_I6/U2_20  ( .A(n970), .B(n589), .CI(
        \position1/sub_226_I6/carry [20]), .CO(
        \position1/sub_226_I6/carry [21]), .S(\position1/N2218 ) );
  ADD32 \position1/sub_226_I7/U2_3  ( .A(n961), .B(n36), .CI(
        \position1/sub_226_I7/carry [3]), .CO(\position1/sub_226_I7/carry [4]), 
        .S(\position1/N2253 ) );
  ADD32 \position1/sub_226_I7/U2_4  ( .A(n960), .B(n245), .CI(
        \position1/sub_226_I7/carry [4]), .CO(\position1/sub_226_I7/carry [5]), 
        .S(\position1/N2254 ) );
  ADD32 \position1/sub_226_I7/U2_5  ( .A(n959), .B(n274), .CI(
        \position1/sub_226_I7/carry [5]), .CO(\position1/sub_226_I7/carry [6]), 
        .S(\position1/N2255 ) );
  ADD32 \position1/sub_226_I7/U2_6  ( .A(n958), .B(n41), .CI(
        \position1/sub_226_I7/carry [6]), .CO(\position1/sub_226_I7/carry [7]), 
        .S(\position1/N2256 ) );
  ADD32 \position1/sub_226_I7/U2_7  ( .A(n957), .B(n278), .CI(
        \position1/sub_226_I7/carry [7]), .CO(\position1/sub_226_I7/carry [8]), 
        .S(\position1/N2257 ) );
  ADD32 \position1/sub_226_I7/U2_8  ( .A(n956), .B(n45), .CI(
        \position1/sub_226_I7/carry [8]), .CO(\position1/sub_226_I7/carry [9]), 
        .S(\position1/N2258 ) );
  ADD32 \position1/sub_226_I7/U2_9  ( .A(n955), .B(n282), .CI(
        \position1/sub_226_I7/carry [9]), .CO(\position1/sub_226_I7/carry [10]), .S(\position1/N2259 ) );
  ADD32 \position1/sub_226_I7/U2_10  ( .A(n954), .B(n40), .CI(
        \position1/sub_226_I7/carry [10]), .CO(
        \position1/sub_226_I7/carry [11]), .S(\position1/N2260 ) );
  ADD32 \position1/sub_226_I7/U2_11  ( .A(n953), .B(n286), .CI(
        \position1/sub_226_I7/carry [11]), .CO(
        \position1/sub_226_I7/carry [12]), .S(\position1/N2261 ) );
  ADD32 \position1/sub_226_I7/U2_12  ( .A(n952), .B(n46), .CI(
        \position1/sub_226_I7/carry [12]), .CO(
        \position1/sub_226_I7/carry [13]), .S(\position1/N2262 ) );
  ADD32 \position1/sub_226_I7/U2_13  ( .A(n951), .B(n261), .CI(
        \position1/sub_226_I7/carry [13]), .CO(
        \position1/sub_226_I7/carry [14]), .S(\position1/N2263 ) );
  ADD32 \position1/sub_226_I7/U2_14  ( .A(n950), .B(n43), .CI(
        \position1/sub_226_I7/carry [14]), .CO(
        \position1/sub_226_I7/carry [15]), .S(\position1/N2264 ) );
  ADD32 \position1/sub_226_I7/U2_15  ( .A(n949), .B(n265), .CI(
        \position1/sub_226_I7/carry [15]), .CO(
        \position1/sub_226_I7/carry [16]), .S(\position1/N2265 ) );
  ADD32 \position1/sub_226_I7/U2_16  ( .A(n948), .B(n42), .CI(
        \position1/sub_226_I7/carry [16]), .CO(
        \position1/sub_226_I7/carry [17]), .S(\position1/N2266 ) );
  ADD32 \position1/sub_226_I7/U2_17  ( .A(n947), .B(n269), .CI(
        \position1/sub_226_I7/carry [17]), .CO(
        \position1/sub_226_I7/carry [18]), .S(\position1/N2267 ) );
  ADD32 \position1/sub_226_I7/U2_18  ( .A(n946), .B(n300), .CI(
        \position1/sub_226_I7/carry [18]), .CO(
        \position1/sub_226_I7/carry [19]), .S(\position1/N2268 ) );
  ADD32 \position1/sub_226_I7/U2_19  ( .A(n945), .B(n590), .CI(
        \position1/sub_226_I7/carry [19]), .CO(
        \position1/sub_226_I7/carry [20]), .S(\position1/N2269 ) );
  ADD32 \position1/sub_226_I8/U2_2  ( .A(n936), .B(n628), .CI(
        \position1/sub_226_I8/carry [2]), .CO(\position1/sub_226_I8/carry [3]), 
        .S(\position1/N2304 ) );
  ADD32 \position1/sub_226_I8/U2_3  ( .A(n934), .B(n272), .CI(
        \position1/sub_226_I8/carry [3]), .CO(\position1/sub_226_I8/carry [4]), 
        .S(\position1/N2305 ) );
  ADD32 \position1/sub_226_I8/U2_4  ( .A(n933), .B(n246), .CI(
        \position1/sub_226_I8/carry [4]), .CO(\position1/sub_226_I8/carry [5]), 
        .S(\position1/N2306 ) );
  ADD32 \position1/sub_226_I8/U2_5  ( .A(n931), .B(n41), .CI(
        \position1/sub_226_I8/carry [5]), .CO(\position1/sub_226_I8/carry [6]), 
        .S(\position1/N2307 ) );
  ADD32 \position1/sub_226_I8/U2_6  ( .A(n930), .B(n250), .CI(
        \position1/sub_226_I8/carry [6]), .CO(\position1/sub_226_I8/carry [7]), 
        .S(\position1/N2308 ) );
  ADD32 \position1/sub_226_I8/U2_7  ( .A(n928), .B(n45), .CI(
        \position1/sub_226_I8/carry [7]), .CO(\position1/sub_226_I8/carry [8]), 
        .S(\position1/N2309 ) );
  ADD32 \position1/sub_226_I8/U2_8  ( .A(n927), .B(n254), .CI(
        \position1/sub_226_I8/carry [8]), .CO(\position1/sub_226_I8/carry [9]), 
        .S(\position1/N2310 ) );
  ADD32 \position1/sub_226_I8/U2_9  ( .A(n925), .B(n40), .CI(
        \position1/sub_226_I8/carry [9]), .CO(\position1/sub_226_I8/carry [10]), .S(\position1/N2311 ) );
  ADD32 \position1/sub_226_I8/U2_10  ( .A(n924), .B(n286), .CI(
        \position1/sub_226_I8/carry [10]), .CO(
        \position1/sub_226_I8/carry [11]), .S(\position1/N2312 ) );
  ADD32 \position1/sub_226_I8/U2_11  ( .A(n923), .B(n46), .CI(
        \position1/sub_226_I8/carry [11]), .CO(
        \position1/sub_226_I8/carry [12]), .S(\position1/N2313 ) );
  ADD32 \position1/sub_226_I8/U2_12  ( .A(n921), .B(n290), .CI(
        \position1/sub_226_I8/carry [12]), .CO(
        \position1/sub_226_I8/carry [13]), .S(\position1/N2314 ) );
  ADD32 \position1/sub_226_I8/U2_13  ( .A(n919), .B(n43), .CI(
        \position1/sub_226_I8/carry [13]), .CO(
        \position1/sub_226_I8/carry [14]), .S(\position1/N2315 ) );
  ADD32 \position1/sub_226_I8/U2_14  ( .A(n918), .B(n294), .CI(
        \position1/sub_226_I8/carry [14]), .CO(
        \position1/sub_226_I8/carry [15]), .S(\position1/N2316 ) );
  ADD32 \position1/sub_226_I8/U2_15  ( .A(n916), .B(n42), .CI(
        \position1/sub_226_I8/carry [15]), .CO(
        \position1/sub_226_I8/carry [16]), .S(\position1/N2317 ) );
  ADD32 \position1/sub_226_I8/U2_16  ( .A(n915), .B(n298), .CI(
        \position1/sub_226_I8/carry [16]), .CO(
        \position1/sub_226_I8/carry [17]), .S(\position1/N2318 ) );
  ADD32 \position1/sub_226_I8/U2_17  ( .A(n914), .B(n44), .CI(
        \position1/sub_226_I8/carry [17]), .CO(
        \position1/sub_226_I8/carry [18]), .S(\position1/N2319 ) );
  ADD32 \position1/sub_226_I8/U2_18  ( .A(n913), .B(n590), .CI(
        \position1/sub_226_I8/carry [18]), .CO(
        \position1/sub_226_I8/carry [19]), .S(\position1/N2320 ) );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_1  ( .A(\position1/x_sum [1]), 
        .B(n835), .CI(\position1/dp_cluster_0/add_196_aco/carry [1]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [2]), .S(\position1/N1178 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_2  ( .A(\position1/x_sum [2]), 
        .B(n855), .CI(\position1/dp_cluster_0/add_196_aco/carry [2]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [3]), .S(\position1/N1179 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_3  ( .A(\position1/x_sum [3]), 
        .B(n857), .CI(\position1/dp_cluster_0/add_196_aco/carry [3]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [4]), .S(\position1/N1180 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_4  ( .A(\position1/x_sum [4]), 
        .B(n859), .CI(\position1/dp_cluster_0/add_196_aco/carry [4]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [5]), .S(\position1/N1181 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_5  ( .A(\position1/x_sum [5]), 
        .B(n861), .CI(\position1/dp_cluster_0/add_196_aco/carry [5]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [6]), .S(\position1/N1182 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_6  ( .A(\position1/x_sum [6]), 
        .B(n863), .CI(\position1/dp_cluster_0/add_196_aco/carry [6]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [7]), .S(\position1/N1183 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_7  ( .A(\position1/x_sum [7]), 
        .B(n866), .CI(\position1/dp_cluster_0/add_196_aco/carry [7]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [8]), .S(\position1/N1184 )
         );
  ADD32 \position1/dp_cluster_0/add_196_aco/U1_8  ( .A(\position1/x_sum [8]), 
        .B(n868), .CI(\position1/dp_cluster_0/add_196_aco/carry [8]), .CO(
        \position1/dp_cluster_0/add_196_aco/carry [9]), .S(\position1/N1185 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_1  ( .A(\position1/y_sum [1]), 
        .B(n808), .CI(\position1/dp_cluster_1/add_197_aco/carry [1]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [2]), .S(\position1/N1203 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_2  ( .A(\position1/y_sum [2]), 
        .B(n804), .CI(\position1/dp_cluster_1/add_197_aco/carry [2]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [3]), .S(\position1/N1204 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_3  ( .A(\position1/y_sum [3]), 
        .B(n800), .CI(\position1/dp_cluster_1/add_197_aco/carry [3]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [4]), .S(\position1/N1205 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_4  ( .A(\position1/y_sum [4]), 
        .B(n796), .CI(\position1/dp_cluster_1/add_197_aco/carry [4]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [5]), .S(\position1/N1206 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_5  ( .A(\position1/y_sum [5]), 
        .B(n792), .CI(\position1/dp_cluster_1/add_197_aco/carry [5]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [6]), .S(\position1/N1207 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_6  ( .A(\position1/y_sum [6]), 
        .B(n788), .CI(\position1/dp_cluster_1/add_197_aco/carry [6]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [7]), .S(\position1/N1208 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_7  ( .A(\position1/y_sum [7]), 
        .B(n784), .CI(\position1/dp_cluster_1/add_197_aco/carry [7]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [8]), .S(\position1/N1209 )
         );
  ADD32 \position1/dp_cluster_1/add_197_aco/U1_8  ( .A(\position1/y_sum [8]), 
        .B(n778), .CI(\position1/dp_cluster_1/add_197_aco/carry [8]), .CO(
        \position1/dp_cluster_1/add_197_aco/carry [9]), .S(\position1/N1210 )
         );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_2  ( .A(
        \position1/N357 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [2]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [3]), .S(
        \position1/N981 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_3  ( .A(
        \position1/N358 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [3]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [4]), .S(
        \position1/N982 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_4  ( .A(
        \position1/N359 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [4]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [5]), .S(
        \position1/N983 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_5  ( .A(
        \position1/N360 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [5]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [6]), .S(
        \position1/N984 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_6  ( .A(
        \position1/N361 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [6]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [7]), .S(
        \position1/N985 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_7  ( .A(
        \position1/N362 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [7]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [8]), .S(
        \position1/N986 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_8  ( .A(
        \position1/N363 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [8]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [9]), .S(
        \position1/N987 ) );
  ADD32 \position1/dp_cluster_2/add_0_root_add_189_3/U1_9  ( .A(
        \position1/N364 ), .B(\position1/dp_cluster_6/N389 ), .CI(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [9]), .CO(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [10]), .S(
        \position1/N988 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_2  ( .A(
        \position1/N282 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [2]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [2]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [3]), .S(
        \position1/N906 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_3  ( .A(
        \position1/N283 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [3]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [3]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [4]), .S(
        \position1/N907 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_4  ( .A(
        \position1/N284 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [4]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [4]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [5]), .S(
        \position1/N908 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_5  ( .A(
        \position1/N285 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [5]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [5]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [6]), .S(
        \position1/N909 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_6  ( .A(
        \position1/N286 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [6]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [6]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [7]), .S(
        \position1/N910 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_7  ( .A(
        \position1/N287 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [7]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [7]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [8]), .S(
        \position1/N911 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_8  ( .A(
        \position1/N288 ), .B(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [8]), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [8]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [9]), .S(
        \position1/N912 ) );
  ADD32 \position1/dp_cluster_3/add_0_root_add_188_3/U1_9  ( .A(
        \position1/N289 ), .B(\position1/dp_cluster_7/N314 ), .CI(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [9]), .CO(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [10]), .S(
        \position1/N913 ) );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_1  ( .A(\position1/x_sum [1]), 
        .B(n834), .CI(\position1/dp_cluster_4/add_178_aco/carry [1]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [2]), .S(\position1/N608 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_2  ( .A(\position1/x_sum [2]), 
        .B(n854), .CI(\position1/dp_cluster_4/add_178_aco/carry [2]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [3]), .S(\position1/N609 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_3  ( .A(\position1/x_sum [3]), 
        .B(n856), .CI(\position1/dp_cluster_4/add_178_aco/carry [3]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [4]), .S(\position1/N610 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_4  ( .A(\position1/x_sum [4]), 
        .B(n858), .CI(\position1/dp_cluster_4/add_178_aco/carry [4]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [5]), .S(\position1/N611 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_5  ( .A(\position1/x_sum [5]), 
        .B(n860), .CI(\position1/dp_cluster_4/add_178_aco/carry [5]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [6]), .S(\position1/N612 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_6  ( .A(\position1/x_sum [6]), 
        .B(n862), .CI(\position1/dp_cluster_4/add_178_aco/carry [6]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [7]), .S(\position1/N613 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_7  ( .A(\position1/x_sum [7]), 
        .B(n865), .CI(\position1/dp_cluster_4/add_178_aco/carry [7]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [8]), .S(\position1/N614 )
         );
  ADD32 \position1/dp_cluster_4/add_178_aco/U1_8  ( .A(\position1/x_sum [8]), 
        .B(n867), .CI(\position1/dp_cluster_4/add_178_aco/carry [8]), .CO(
        \position1/dp_cluster_4/add_178_aco/carry [9]), .S(\position1/N615 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_1  ( .A(\position1/y_sum [1]), 
        .B(n807), .CI(\position1/dp_cluster_5/add_179_aco/carry [1]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [2]), .S(\position1/N633 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_2  ( .A(\position1/y_sum [2]), 
        .B(n803), .CI(\position1/dp_cluster_5/add_179_aco/carry [2]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [3]), .S(\position1/N634 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_3  ( .A(\position1/y_sum [3]), 
        .B(n799), .CI(\position1/dp_cluster_5/add_179_aco/carry [3]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [4]), .S(\position1/N635 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_4  ( .A(\position1/y_sum [4]), 
        .B(n795), .CI(\position1/dp_cluster_5/add_179_aco/carry [4]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [5]), .S(\position1/N636 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_5  ( .A(\position1/y_sum [5]), 
        .B(n791), .CI(\position1/dp_cluster_5/add_179_aco/carry [5]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [6]), .S(\position1/N637 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_6  ( .A(\position1/y_sum [6]), 
        .B(n787), .CI(\position1/dp_cluster_5/add_179_aco/carry [6]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [7]), .S(\position1/N638 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_7  ( .A(\position1/y_sum [7]), 
        .B(n783), .CI(\position1/dp_cluster_5/add_179_aco/carry [7]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [8]), .S(\position1/N639 )
         );
  ADD32 \position1/dp_cluster_5/add_179_aco/U1_8  ( .A(\position1/y_sum [8]), 
        .B(n777), .CI(\position1/dp_cluster_5/add_179_aco/carry [8]), .CO(
        \position1/dp_cluster_5/add_179_aco/carry [9]), .S(\position1/N640 )
         );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_2  ( .A(
        \position1/N357 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [2]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [3]), .S(
        \position1/N407 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_3  ( .A(
        \position1/N358 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [3]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [4]), .S(
        \position1/N408 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_4  ( .A(
        \position1/N359 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [4]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [5]), .S(
        \position1/N409 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_5  ( .A(
        \position1/N360 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [5]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [6]), .S(
        \position1/N410 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_6  ( .A(
        \position1/N361 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [6]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [7]), .S(
        \position1/N411 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_7  ( .A(
        \position1/N362 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [7]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [8]), .S(
        \position1/N412 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_8  ( .A(
        \position1/N363 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [8]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [9]), .S(
        \position1/N413 ) );
  ADD32 \position1/dp_cluster_6/add_0_root_add_171_3/U1_9  ( .A(
        \position1/N364 ), .B(\position1/dp_cluster_6/N389 ), .CI(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [9]), .CO(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [10]), .S(
        \position1/N414 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_2  ( .A(
        \position1/N282 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [2]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [2]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [3]), .S(
        \position1/N332 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_3  ( .A(
        \position1/N283 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [3]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [3]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [4]), .S(
        \position1/N333 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_4  ( .A(
        \position1/N284 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [4]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [4]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [5]), .S(
        \position1/N334 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_5  ( .A(
        \position1/N285 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [5]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [5]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [6]), .S(
        \position1/N335 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_6  ( .A(
        \position1/N286 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [6]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [6]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [7]), .S(
        \position1/N336 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_7  ( .A(
        \position1/N287 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [7]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [7]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [8]), .S(
        \position1/N337 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_8  ( .A(
        \position1/N288 ), .B(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [8]), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [8]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [9]), .S(
        \position1/N338 ) );
  ADD32 \position1/dp_cluster_7/add_0_root_add_170_3/U1_9  ( .A(
        \position1/N289 ), .B(\position1/dp_cluster_7/N314 ), .CI(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [9]), .CO(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [10]), .S(
        \position1/N339 ) );
  ADD22 \gensync1/add_39/U1_1_1  ( .A(\gensync1/N182 ), .B(\gensync1/N74 ), 
        .CO(\gensync1/add_39/carry [2]), .S(\gensync1/N13 ) );
  ADD22 \gensync1/add_39/U1_1_2  ( .A(\gensync1/N181 ), .B(
        \gensync1/add_39/carry [2]), .CO(\gensync1/add_39/carry [3]), .S(
        \gensync1/N14 ) );
  ADD22 \gensync1/add_39/U1_1_3  ( .A(\gensync1/N180 ), .B(
        \gensync1/add_39/carry [3]), .CO(\gensync1/add_39/carry [4]), .S(
        \gensync1/N15 ) );
  ADD22 \gensync1/add_39/U1_1_4  ( .A(\gensync1/N179 ), .B(
        \gensync1/add_39/carry [4]), .CO(\gensync1/add_39/carry [5]), .S(
        \gensync1/N16 ) );
  ADD22 \gensync1/add_39/U1_1_5  ( .A(\gensync1/N178 ), .B(
        \gensync1/add_39/carry [5]), .CO(\gensync1/add_39/carry [6]), .S(
        \gensync1/N17 ) );
  ADD22 \gensync1/add_39/U1_1_6  ( .A(\gensync1/N177 ), .B(
        \gensync1/add_39/carry [6]), .CO(\gensync1/add_39/carry [7]), .S(
        \gensync1/N18 ) );
  ADD22 \gensync1/add_39/U1_1_7  ( .A(\gensync1/N176 ), .B(
        \gensync1/add_39/carry [7]), .CO(\gensync1/add_39/carry [8]), .S(
        \gensync1/N19 ) );
  ADD22 \gensync1/add_39/U1_1_8  ( .A(\gensync1/N175 ), .B(
        \gensync1/add_39/carry [8]), .CO(\gensync1/add_39/carry [9]), .S(
        \gensync1/N20 ) );
  ADD22 \gensync1/add_45/U1_1_1  ( .A(\gensync1/N172 ), .B(\gensync1/N173 ), 
        .CO(\gensync1/add_45/carry [2]), .S(\gensync1/N47 ) );
  ADD22 \gensync1/add_45/U1_1_2  ( .A(\gensync1/N171 ), .B(
        \gensync1/add_45/carry [2]), .CO(\gensync1/add_45/carry [3]), .S(
        \gensync1/N48 ) );
  ADD22 \gensync1/add_45/U1_1_3  ( .A(\gensync1/N170 ), .B(
        \gensync1/add_45/carry [3]), .CO(\gensync1/add_45/carry [4]), .S(
        \gensync1/N49 ) );
  ADD22 \gensync1/add_45/U1_1_4  ( .A(\gensync1/N169 ), .B(
        \gensync1/add_45/carry [4]), .CO(\gensync1/add_45/carry [5]), .S(
        \gensync1/N50 ) );
  ADD22 \gensync1/add_45/U1_1_5  ( .A(\gensync1/N168 ), .B(
        \gensync1/add_45/carry [5]), .CO(\gensync1/add_45/carry [6]), .S(
        \gensync1/N51 ) );
  ADD22 \gensync1/add_45/U1_1_6  ( .A(\gensync1/N167 ), .B(
        \gensync1/add_45/carry [6]), .CO(\gensync1/add_45/carry [7]), .S(
        \gensync1/N52 ) );
  ADD22 \gensync1/add_45/U1_1_7  ( .A(\gensync1/N166 ), .B(
        \gensync1/add_45/carry [7]), .CO(\gensync1/add_45/carry [8]), .S(
        \gensync1/N53 ) );
  ADD22 \gensync1/add_45/U1_1_8  ( .A(\gensync1/N165 ), .B(
        \gensync1/add_45/carry [8]), .CO(\gensync1/add_45/carry [9]), .S(
        \gensync1/N54 ) );
  DF3 \gensync1/VSYNC_reg  ( .D(n815), .C(CLK_top), .Q(VSYNC_top) );
  DF3 \gensync1/HSYNC_reg  ( .D(n872), .C(CLK_top), .Q(HSYNC_top) );
  DF3 \gensync1/comptX_reg[1]  ( .D(\gensync1/N23 ), .C(CLK_top), .Q(
        \gensync1/N182 ), .QN(n10) );
  DF3 \gensync1/comptX_reg[2]  ( .D(\gensync1/N24 ), .C(CLK_top), .Q(
        \gensync1/N181 ), .QN(n4) );
  DF3 \gensync1/comptX_reg[3]  ( .D(\gensync1/N25 ), .C(CLK_top), .Q(
        \gensync1/N180 ), .QN(n12) );
  DF3 \gensync1/comptX_reg[4]  ( .D(\gensync1/N26 ), .C(CLK_top), .Q(
        \gensync1/N179 ), .QN(n7) );
  DF3 \gensync1/comptX_reg[5]  ( .D(\gensync1/N27 ), .C(CLK_top), .Q(
        \gensync1/N178 ), .QN(n14) );
  DF3 \gensync1/comptX_reg[6]  ( .D(\gensync1/N28 ), .C(CLK_top), .Q(
        \gensync1/N177 ), .QN(n6) );
  DF3 \gensync1/comptX_reg[7]  ( .D(\gensync1/N29 ), .C(CLK_top), .Q(
        \gensync1/N176 ), .QN(n15) );
  DF3 \gensync1/comptX_reg[8]  ( .D(\gensync1/N30 ), .C(CLK_top), .Q(
        \gensync1/N175 ) );
  DF3 \gensync1/comptX_reg[9]  ( .D(\gensync1/N31 ), .C(CLK_top), .Q(
        \gensync1/N174 ) );
  DF3 \gensync1/comptX_reg[0]  ( .D(\gensync1/N22 ), .C(CLK_top), .Q(
        \gensync1/N74 ), .QN(n1) );
  DF3 \image_process1/state_reg  ( .D(reset_top), .C(CLK_top), .Q(
        \image_process1/state ), .QN(\image_process1/n27 ) );
  DF3 \image_process1/bi_reg[0]  ( .D(n749), .C(CLK_top), .Q(
        \image_process1/bi [0]) );
  DF3 \image_process1/bi_reg[1]  ( .D(n748), .C(CLK_top), .Q(
        \image_process1/bi [1]) );
  DF3 \image_process1/bi_reg[2]  ( .D(n747), .C(CLK_top), .QN(
        \image_process1/n25 ) );
  DF3 \image_process1/bi_reg[3]  ( .D(n746), .C(CLK_top), .Q(
        \image_process1/bi [3]) );
  DF3 \image_process1/bi_reg[4]  ( .D(n745), .C(CLK_top), .Q(
        \image_process1/bi [4]) );
  DF3 \image_process1/bi_reg[5]  ( .D(n744), .C(CLK_top), .Q(
        \image_process1/bi [5]) );
  DF3 \image_process1/bi_reg[6]  ( .D(n743), .C(CLK_top), .Q(
        \image_process1/bi [6]) );
  DF3 \image_process1/bi_reg[7]  ( .D(n742), .C(CLK_top), .Q(
        \image_process1/bi [7]) );
  DF3 \image_process1/gi_reg[0]  ( .D(n757), .C(CLK_top), .Q(
        \image_process1/gi [0]) );
  DF3 \image_process1/gi_reg[1]  ( .D(n756), .C(CLK_top), .Q(
        \image_process1/gi [1]) );
  DF3 \image_process1/gi_reg[2]  ( .D(n755), .C(CLK_top), .Q(
        \image_process1/gi [2]) );
  DF3 \image_process1/gi_reg[3]  ( .D(n754), .C(CLK_top), .Q(
        \image_process1/gi [3]) );
  DF3 \image_process1/gi_reg[4]  ( .D(n753), .C(CLK_top), .Q(
        \image_process1/gi [4]), .QN(n5) );
  DF3 \image_process1/gi_reg[5]  ( .D(n752), .C(CLK_top), .Q(
        \image_process1/gi [5]), .QN(n33) );
  DF3 \image_process1/gi_reg[6]  ( .D(n751), .C(CLK_top), .Q(
        \image_process1/gi [6]) );
  DF3 \image_process1/gi_reg[7]  ( .D(n750), .C(CLK_top), .Q(
        \image_process1/gi [7]) );
  DF3 \image_process1/ri_reg[0]  ( .D(n765), .C(CLK_top), .Q(
        \image_process1/ri [0]) );
  DF3 \image_process1/ri_reg[1]  ( .D(n764), .C(CLK_top), .Q(
        \image_process1/ri [1]) );
  DF3 \image_process1/ri_reg[2]  ( .D(n763), .C(CLK_top), .QN(
        \image_process1/n13 ) );
  DF3 \image_process1/ri_reg[3]  ( .D(n762), .C(CLK_top), .Q(
        \image_process1/ri [3]) );
  DF3 \image_process1/ri_reg[4]  ( .D(n761), .C(CLK_top), .Q(
        \image_process1/ri [4]) );
  DF3 \image_process1/ri_reg[5]  ( .D(n760), .C(CLK_top), .Q(
        \image_process1/ri [5]) );
  DF3 \image_process1/ri_reg[6]  ( .D(n759), .C(CLK_top), .Q(
        \image_process1/ri [6]) );
  DF3 \image_process1/ri_reg[7]  ( .D(n758), .C(CLK_top), .Q(
        \image_process1/ri [7]) );
  DF3 \position1/b_bout_reg[3]  ( .D(\position1/N100 ), .C(CLK_top), .Q(
        bout_top[3]) );
  DF3 \position1/b_bout_reg[4]  ( .D(\position1/N101 ), .C(CLK_top), .Q(
        bout_top[4]) );
  DF3 \position1/b_bout_reg[5]  ( .D(\position1/N102 ), .C(CLK_top), .Q(
        bout_top[5]) );
  DF3 \position1/b_bout_reg[6]  ( .D(\position1/N103 ), .C(CLK_top), .Q(
        bout_top[6]) );
  DF3 \position1/b_bout_reg[7]  ( .D(\position1/N104 ), .C(CLK_top), .Q(
        bout_top[7]) );
  DF3 \position1/r_bout_reg[0]  ( .D(\position1/N81 ), .C(CLK_top), .Q(
        rout_top[0]) );
  DF3 \position1/r_bout_reg[1]  ( .D(\position1/N82 ), .C(CLK_top), .Q(
        rout_top[1]) );
  DF3 \position1/r_bout_reg[2]  ( .D(\position1/N83 ), .C(CLK_top), .Q(
        rout_top[2]) );
  DF3 \position1/r_bout_reg[3]  ( .D(\position1/N84 ), .C(CLK_top), .Q(
        rout_top[3]) );
  DF3 \position1/r_bout_reg[4]  ( .D(\position1/N85 ), .C(CLK_top), .Q(
        rout_top[4]) );
  DF3 \position1/r_bout_reg[5]  ( .D(\position1/N86 ), .C(CLK_top), .Q(
        rout_top[5]) );
  DF3 \position1/r_bout_reg[6]  ( .D(\position1/N87 ), .C(CLK_top), .Q(
        rout_top[6]) );
  DF3 \position1/r_bout_reg[7]  ( .D(\position1/N88 ), .C(CLK_top), .Q(
        rout_top[7]) );
  DF3 \position1/b_bout_reg[0]  ( .D(\position1/N97 ), .C(CLK_top), .Q(
        bout_top[0]) );
  DF3 \position1/b_bout_reg[1]  ( .D(\position1/N98 ), .C(CLK_top), .Q(
        bout_top[1]) );
  DF3 \position1/b_bout_reg[2]  ( .D(\position1/N99 ), .C(CLK_top), .Q(
        bout_top[2]) );
  DF3 \position1/g_bout_reg[1]  ( .D(n713), .C(CLK_top), .Q(gout_top[1]) );
  DF3 \position1/g_bout_reg[3]  ( .D(n714), .C(CLK_top), .Q(gout_top[3]) );
  DF3 \position1/g_bout_reg[7]  ( .D(n715), .C(CLK_top), .Q(gout_top[7]) );
  DF3 \position1/g_bout_reg[0]  ( .D(\position1/N89 ), .C(CLK_top), .Q(
        gout_top[0]) );
  DF3 \position1/g_bout_reg[2]  ( .D(\position1/N91 ), .C(CLK_top), .Q(
        gout_top[2]) );
  DF3 \position1/g_bout_reg[4]  ( .D(\position1/N93 ), .C(CLK_top), .Q(
        gout_top[4]) );
  DF3 \position1/g_bout_reg[5]  ( .D(\position1/N94 ), .C(CLK_top), .Q(
        gout_top[5]) );
  DF3 \position1/g_bout_reg[6]  ( .D(\position1/N95 ), .C(CLK_top), .Q(
        gout_top[6]) );
  DF3 \position1/y_bar_reg[0]  ( .D(n683), .C(CLK_top), .Q(Y_barycentre_top[0]) );
  DLPQ3 \position1/quot_y_reg[0]  ( .SN(\position1/n283 ), .D(
        \position1/N2363 ), .GN(n1358), .Q(\position1/quot_y [0]) );
  DF3 \position1/y_bar_reg[1]  ( .D(n684), .C(CLK_top), .Q(Y_barycentre_top[1]), .QN(n23) );
  DLPQ3 \position1/quot_y_reg[1]  ( .SN(\position1/n283 ), .D(
        \position1/N2364 ), .GN(n1358), .Q(\position1/quot_y [1]) );
  DF3 \position1/y_bar_reg[2]  ( .D(n685), .C(CLK_top), .Q(Y_barycentre_top[2]), .QN(n21) );
  DLPQ3 \position1/quot_y_reg[2]  ( .SN(\position1/n283 ), .D(
        \position1/N2365 ), .GN(n1358), .Q(\position1/quot_y [2]) );
  DF3 \position1/y_bar_reg[3]  ( .D(n686), .C(CLK_top), .Q(Y_barycentre_top[3]), .QN(n24) );
  DLPQ3 \position1/quot_y_reg[3]  ( .SN(\position1/n283 ), .D(
        \position1/N2366 ), .GN(n1358), .Q(\position1/quot_y [3]) );
  DF3 \position1/y_bar_reg[4]  ( .D(n687), .C(CLK_top), .Q(Y_barycentre_top[4]), .QN(n26) );
  DLPQ3 \position1/quot_y_reg[4]  ( .SN(\position1/n283 ), .D(
        \position1/N2367 ), .GN(n1358), .Q(\position1/quot_y [4]) );
  DF3 \position1/y_bar_reg[5]  ( .D(n688), .C(CLK_top), .Q(Y_barycentre_top[5]), .QN(n28) );
  DLPQ3 \position1/quot_y_reg[5]  ( .SN(\position1/n283 ), .D(
        \position1/N2368 ), .GN(n1358), .Q(\position1/quot_y [5]) );
  DF3 \position1/y_bar_reg[6]  ( .D(n689), .C(CLK_top), .Q(Y_barycentre_top[6]), .QN(n31) );
  DLPQ3 \position1/quot_y_reg[6]  ( .SN(\position1/n283 ), .D(
        \position1/N2369 ), .GN(n1358), .Q(\position1/quot_y [6]) );
  DF3 \position1/y_bar_reg[7]  ( .D(n690), .C(CLK_top), .Q(Y_barycentre_top[7]), .QN(n32) );
  DLPQ3 \position1/quot_y_reg[7]  ( .SN(\position1/n283 ), .D(
        \position1/N2370 ), .GN(n1358), .Q(\position1/quot_y [7]) );
  DF3 \position1/y_bar_reg[8]  ( .D(n691), .C(CLK_top), .Q(Y_barycentre_top[8]), .QN(n30) );
  DLPQ3 \position1/quot_y_reg[8]  ( .SN(\position1/n283 ), .D(
        \position1/N2371 ), .GN(n1358), .Q(\position1/quot_y [8]) );
  DF3 \position1/x_bar_reg[0]  ( .D(n674), .C(CLK_top), .Q(X_barycentre_top[0]) );
  DLPQ3 \position1/quot_x_reg[0]  ( .SN(\position1/n283 ), .D(
        \position1/N2354 ), .GN(n1358), .Q(\position1/quot_x [0]) );
  DF3 \position1/x_bar_reg[1]  ( .D(n675), .C(CLK_top), .Q(X_barycentre_top[1]), .QN(n17) );
  DLPQ3 \position1/quot_x_reg[1]  ( .SN(\position1/n283 ), .D(
        \position1/N2355 ), .GN(n1358), .Q(\position1/quot_x [1]) );
  DF3 \position1/x_bar_reg[2]  ( .D(n676), .C(CLK_top), .Q(X_barycentre_top[2]), .QN(n16) );
  DLPQ3 \position1/quot_x_reg[2]  ( .SN(\position1/n283 ), .D(
        \position1/N2356 ), .GN(n1358), .Q(\position1/quot_x [2]) );
  DF3 \position1/x_bar_reg[3]  ( .D(n677), .C(CLK_top), .Q(X_barycentre_top[3]), .QN(n19) );
  DLPQ3 \position1/quot_x_reg[3]  ( .SN(\position1/n283 ), .D(
        \position1/N2357 ), .GN(n1358), .Q(\position1/quot_x [3]) );
  DF3 \position1/x_bar_reg[4]  ( .D(n678), .C(CLK_top), .Q(X_barycentre_top[4]), .QN(n20) );
  DLPQ3 \position1/quot_x_reg[4]  ( .SN(\position1/n283 ), .D(
        \position1/N2358 ), .GN(n1358), .Q(\position1/quot_x [4]) );
  DF3 \position1/x_bar_reg[5]  ( .D(n679), .C(CLK_top), .Q(X_barycentre_top[5]), .QN(n22) );
  DLPQ3 \position1/quot_x_reg[5]  ( .SN(\position1/n283 ), .D(
        \position1/N2359 ), .GN(n1358), .Q(\position1/quot_x [5]) );
  DF3 \position1/x_bar_reg[6]  ( .D(n680), .C(CLK_top), .Q(X_barycentre_top[6]), .QN(n25) );
  DLPQ3 \position1/quot_x_reg[6]  ( .SN(\position1/n283 ), .D(
        \position1/N2360 ), .GN(n1358), .Q(\position1/quot_x [6]) );
  DF3 \position1/x_bar_reg[7]  ( .D(n681), .C(CLK_top), .Q(X_barycentre_top[7]), .QN(n27) );
  DLPQ3 \position1/quot_x_reg[7]  ( .SN(\position1/n283 ), .D(
        \position1/N2361 ), .GN(n1358), .Q(\position1/quot_x [7]) );
  DF3 \position1/x_bar_reg[8]  ( .D(n682), .C(CLK_top), .Q(X_barycentre_top[8]), .QN(n29) );
  DLPQ3 \position1/quot_x_reg[8]  ( .SN(\position1/n283 ), .D(
        \position1/N2362 ), .GN(n1358), .Q(\position1/quot_x [8]) );
  DF3 \position1/count_reg[15]  ( .D(n670), .C(CLK_top), .Q(\position1/N2446 ), 
        .QN(n67) );
  DF3 \position1/count_reg[14]  ( .D(n669), .C(CLK_top), .Q(\position1/N2447 ), 
        .QN(n42) );
  DF3 \position1/count_reg[13]  ( .D(n668), .C(CLK_top), .Q(\position1/N2448 ), 
        .QN(n39) );
  DF3 \position1/count_reg[12]  ( .D(n667), .C(CLK_top), .Q(\position1/N2449 ), 
        .QN(n43) );
  DF3 \position1/count_reg[11]  ( .D(n666), .C(CLK_top), .Q(\position1/N2450 ), 
        .QN(n38) );
  DF3 \position1/count_reg[10]  ( .D(n665), .C(CLK_top), .Q(\position1/N2451 ), 
        .QN(n46) );
  DF3 \position1/count_reg[9]  ( .D(n664), .C(CLK_top), .Q(\position1/N2452 ), 
        .QN(n35) );
  DF3 \position1/count_reg[8]  ( .D(n663), .C(CLK_top), .Q(\position1/N2453 ), 
        .QN(n40) );
  DF3 \position1/count_reg[7]  ( .D(n662), .C(CLK_top), .Q(\position1/N2454 ), 
        .QN(n100) );
  DF3 \position1/count_reg[6]  ( .D(n661), .C(CLK_top), .Q(\position1/N2455 ), 
        .QN(n45) );
  DF3 \position1/count_reg[5]  ( .D(n660), .C(CLK_top), .Q(\position1/N2456 ), 
        .QN(n47) );
  DF3 \position1/count_reg[4]  ( .D(n659), .C(CLK_top), .Q(\position1/N2457 ), 
        .QN(n41) );
  DF3 \position1/count_reg[3]  ( .D(n658), .C(CLK_top), .Q(\position1/N2458 ), 
        .QN(n37) );
  DF3 \position1/count_reg[2]  ( .D(n657), .C(CLK_top), .Q(\position1/N2459 ), 
        .QN(n66) );
  DF3 \position1/count_reg[1]  ( .D(n656), .C(CLK_top), .Q(\position1/N2460 ), 
        .QN(n36) );
  DF3 \position1/count_reg[16]  ( .D(n671), .C(CLK_top), .Q(\position1/N2445 ), 
        .QN(n44) );
  DF3 \position1/count_reg[17]  ( .D(n672), .C(CLK_top), .Q(n2), .QN(n101) );
  DF3 \position1/count_reg[0]  ( .D(n655), .C(CLK_top), .Q(\position1/N560 ), 
        .QN(n34) );
  DF3 \position1/x_sum_reg[22]  ( .D(\position1/n1613 ), .C(CLK_top), .Q(
        \position1/x_sum [22]), .QN(n76) );
  DF3 \position1/x_sum_reg[21]  ( .D(\position1/n1614 ), .C(CLK_top), .Q(
        \position1/x_sum [21]), .QN(n60) );
  DF3 \position1/x_sum_reg[20]  ( .D(\position1/n1615 ), .C(CLK_top), .Q(
        \position1/x_sum [20]), .QN(n77) );
  DF3 \position1/x_sum_reg[19]  ( .D(\position1/n1616 ), .C(CLK_top), .Q(
        \position1/x_sum [19]), .QN(n61) );
  DF3 \position1/x_sum_reg[18]  ( .D(\position1/n1617 ), .C(CLK_top), .Q(
        \position1/x_sum [18]), .QN(n78) );
  DF3 \position1/x_sum_reg[17]  ( .D(\position1/n1618 ), .C(CLK_top), .Q(
        \position1/x_sum [17]), .QN(n62) );
  DF3 \position1/x_sum_reg[16]  ( .D(\position1/n1619 ), .C(CLK_top), .Q(
        \position1/x_sum [16]), .QN(n79) );
  DF3 \position1/x_sum_reg[15]  ( .D(\position1/n1620 ), .C(CLK_top), .Q(
        \position1/x_sum [15]), .QN(n63) );
  DF3 \position1/x_sum_reg[14]  ( .D(\position1/n1621 ), .C(CLK_top), .Q(
        \position1/x_sum [14]), .QN(n80) );
  DF3 \position1/x_sum_reg[13]  ( .D(\position1/n1622 ), .C(CLK_top), .Q(
        \position1/x_sum [13]), .QN(n64) );
  DF3 \position1/x_sum_reg[12]  ( .D(\position1/n1623 ), .C(CLK_top), .Q(
        \position1/x_sum [12]), .QN(n81) );
  DF3 \position1/x_sum_reg[11]  ( .D(\position1/n1624 ), .C(CLK_top), .Q(
        \position1/x_sum [11]), .QN(n65) );
  DF3 \position1/x_sum_reg[10]  ( .D(\position1/n1625 ), .C(CLK_top), .Q(
        \position1/x_sum [10]), .QN(n69) );
  DF3 \position1/x_sum_reg[9]  ( .D(\position1/n1626 ), .C(CLK_top), .Q(
        \position1/x_sum [9]), .QN(n51) );
  DF3 \position1/x_sum_reg[8]  ( .D(\position1/n1627 ), .C(CLK_top), .Q(
        \position1/x_sum [8]), .QN(n49) );
  DF3 \position1/x_sum_reg[7]  ( .D(\position1/n1628 ), .C(CLK_top), .Q(
        \position1/x_sum [7]), .QN(n94) );
  DF3 \position1/x_sum_reg[6]  ( .D(\position1/n1629 ), .C(CLK_top), .Q(
        \position1/x_sum [6]), .QN(n87) );
  DF3 \position1/x_sum_reg[5]  ( .D(\position1/n1630 ), .C(CLK_top), .Q(
        \position1/x_sum [5]), .QN(n88) );
  DF3 \position1/x_sum_reg[4]  ( .D(\position1/n1631 ), .C(CLK_top), .Q(
        \position1/x_sum [4]), .QN(n89) );
  DF3 \position1/x_sum_reg[3]  ( .D(\position1/n1632 ), .C(CLK_top), .Q(
        \position1/x_sum [3]), .QN(n95) );
  DF3 \position1/x_sum_reg[2]  ( .D(\position1/n1633 ), .C(CLK_top), .Q(
        \position1/x_sum [2]), .QN(n90) );
  DF3 \position1/x_sum_reg[1]  ( .D(\position1/n1634 ), .C(CLK_top), .Q(
        \position1/x_sum [1]), .QN(n91) );
  DF3 \position1/x_sum_reg[23]  ( .D(\position1/n1612 ), .C(CLK_top), .Q(
        \position1/x_sum [23]), .QN(n59) );
  DF3 \position1/x_sum_reg[24]  ( .D(\position1/n1611 ), .C(CLK_top), .Q(
        \position1/x_sum [24]), .QN(n99) );
  DF3 \position1/x_sum_reg[0]  ( .D(\position1/n1635 ), .C(CLK_top), .Q(
        \position1/N1521 ), .QN(n97) );
  DF3 \position1/y_sum_reg[22]  ( .D(\position1/n1588 ), .C(CLK_top), .Q(
        \position1/y_sum [22]), .QN(n70) );
  DF3 \position1/y_sum_reg[21]  ( .D(\position1/n1589 ), .C(CLK_top), .Q(
        \position1/y_sum [21]), .QN(n53) );
  DF3 \position1/y_sum_reg[20]  ( .D(\position1/n1590 ), .C(CLK_top), .Q(
        \position1/y_sum [20]), .QN(n71) );
  DF3 \position1/y_sum_reg[19]  ( .D(\position1/n1591 ), .C(CLK_top), .Q(
        \position1/y_sum [19]), .QN(n54) );
  DF3 \position1/y_sum_reg[18]  ( .D(\position1/n1592 ), .C(CLK_top), .Q(
        \position1/y_sum [18]), .QN(n72) );
  DF3 \position1/y_sum_reg[17]  ( .D(\position1/n1593 ), .C(CLK_top), .Q(
        \position1/y_sum [17]), .QN(n55) );
  DF3 \position1/y_sum_reg[16]  ( .D(\position1/n1594 ), .C(CLK_top), .Q(
        \position1/y_sum [16]), .QN(n73) );
  DF3 \position1/y_sum_reg[15]  ( .D(\position1/n1595 ), .C(CLK_top), .Q(
        \position1/y_sum [15]), .QN(n56) );
  DF3 \position1/y_sum_reg[14]  ( .D(\position1/n1596 ), .C(CLK_top), .Q(
        \position1/y_sum [14]), .QN(n74) );
  DF3 \position1/y_sum_reg[13]  ( .D(\position1/n1597 ), .C(CLK_top), .Q(
        \position1/y_sum [13]), .QN(n57) );
  DF3 \position1/y_sum_reg[12]  ( .D(\position1/n1598 ), .C(CLK_top), .Q(
        \position1/y_sum [12]), .QN(n75) );
  DF3 \position1/y_sum_reg[11]  ( .D(\position1/n1599 ), .C(CLK_top), .Q(
        \position1/y_sum [11]), .QN(n58) );
  DF3 \position1/y_sum_reg[10]  ( .D(\position1/n1600 ), .C(CLK_top), .Q(
        \position1/y_sum [10]), .QN(n68) );
  DF3 \position1/y_sum_reg[9]  ( .D(\position1/n1601 ), .C(CLK_top), .Q(
        \position1/y_sum [9]), .QN(n50) );
  DF3 \position1/y_sum_reg[8]  ( .D(\position1/n1602 ), .C(CLK_top), .Q(
        \position1/y_sum [8]), .QN(n48) );
  DF3 \position1/y_sum_reg[7]  ( .D(\position1/n1603 ), .C(CLK_top), .Q(
        \position1/y_sum [7]), .QN(n92) );
  DF3 \position1/y_sum_reg[6]  ( .D(\position1/n1604 ), .C(CLK_top), .Q(
        \position1/y_sum [6]), .QN(n82) );
  DF3 \position1/y_sum_reg[5]  ( .D(\position1/n1605 ), .C(CLK_top), .Q(
        \position1/y_sum [5]), .QN(n83) );
  DF3 \position1/y_sum_reg[4]  ( .D(\position1/n1606 ), .C(CLK_top), .Q(
        \position1/y_sum [4]), .QN(n84) );
  DF3 \position1/y_sum_reg[3]  ( .D(\position1/n1607 ), .C(CLK_top), .Q(
        \position1/y_sum [3]), .QN(n93) );
  DF3 \position1/y_sum_reg[2]  ( .D(\position1/n1608 ), .C(CLK_top), .Q(
        \position1/y_sum [2]), .QN(n85) );
  DF3 \position1/y_sum_reg[1]  ( .D(\position1/n1609 ), .C(CLK_top), .Q(
        \position1/y_sum [1]), .QN(n86) );
  DF3 \position1/y_sum_reg[23]  ( .D(\position1/n1587 ), .C(CLK_top), .Q(
        \position1/y_sum [23]), .QN(n52) );
  DF3 \position1/y_sum_reg[24]  ( .D(\position1/n1586 ), .C(CLK_top), .Q(
        \position1/y_sum [24]), .QN(n98) );
  DF3 \position1/y_sum_reg[0]  ( .D(\position1/n1610 ), .C(CLK_top), .Q(
        \position1/N1938 ), .QN(n96) );
  DF3 \position1/count_img_reg[19]  ( .D(n711), .C(CLK_top), .Q(
        \position1/count_img [19]) );
  DF3 \position1/count_img_reg[18]  ( .D(n710), .C(CLK_top), .Q(
        \position1/count_img [18]) );
  DF3 \position1/count_img_reg[17]  ( .D(n709), .C(CLK_top), .Q(
        \position1/count_img [17]) );
  DF3 \position1/count_img_reg[16]  ( .D(n708), .C(CLK_top), .Q(
        \position1/count_img [16]) );
  DF3 \position1/count_img_reg[15]  ( .D(n707), .C(CLK_top), .Q(
        \position1/count_img [15]), .QN(n18) );
  DF3 \position1/count_img_reg[14]  ( .D(n706), .C(CLK_top), .Q(
        \position1/count_img [14]) );
  DF3 \position1/count_img_reg[13]  ( .D(n705), .C(CLK_top), .Q(
        \position1/count_img [13]) );
  DF3 \position1/count_img_reg[12]  ( .D(n704), .C(CLK_top), .Q(
        \position1/count_img [12]) );
  DF3 \position1/count_img_reg[11]  ( .D(n703), .C(CLK_top), .Q(
        \position1/count_img [11]) );
  DF3 \position1/count_img_reg[10]  ( .D(n702), .C(CLK_top), .Q(
        \position1/count_img [10]) );
  DF3 \position1/count_img_reg[9]  ( .D(n701), .C(CLK_top), .Q(
        \position1/count_img [9]) );
  DF3 \position1/count_img_reg[8]  ( .D(n700), .C(CLK_top), .Q(
        \position1/count_img [8]) );
  DF3 \position1/count_img_reg[7]  ( .D(n699), .C(CLK_top), .Q(
        \position1/count_img [7]) );
  DF3 \position1/count_img_reg[6]  ( .D(n698), .C(CLK_top), .Q(
        \position1/count_img [6]) );
  DF3 \position1/count_img_reg[5]  ( .D(n697), .C(CLK_top), .Q(
        \position1/count_img [5]) );
  DF3 \position1/count_img_reg[4]  ( .D(n696), .C(CLK_top), .Q(
        \position1/count_img [4]) );
  DF3 \position1/count_img_reg[3]  ( .D(n695), .C(CLK_top), .Q(
        \position1/count_img [3]) );
  DF3 \position1/count_img_reg[2]  ( .D(n694), .C(CLK_top), .Q(
        \position1/count_img [2]) );
  DF3 \position1/count_img_reg[1]  ( .D(n693), .C(CLK_top), .Q(
        \position1/count_img [1]) );
  DF3 \position1/state_reg[1]  ( .D(n484), .C(CLK_top), .Q(
        \position1/state [1]), .QN(\position1/n344 ) );
  DF3 \position1/state_reg[0]  ( .D(\position1/N193 ), .C(CLK_top), .Q(
        \position1/state [0]) );
  DF3 \position1/count_img_reg[0]  ( .D(n692), .C(CLK_top), .Q(
        \position1/count_img [0]), .QN(\position1/n802 ) );
  DF3 \position1/bi_reg[0]  ( .D(n723), .C(CLK_top), .QN(\position1/n370 ) );
  DF3 \position1/bi_reg[1]  ( .D(n722), .C(CLK_top), .QN(\position1/n369 ) );
  DF3 \position1/bi_reg[2]  ( .D(n721), .C(CLK_top), .QN(\position1/n368 ) );
  DF3 \position1/bi_reg[3]  ( .D(n720), .C(CLK_top), .QN(\position1/n367 ) );
  DF3 \position1/bi_reg[4]  ( .D(n719), .C(CLK_top), .QN(\position1/n366 ) );
  DF3 \position1/bi_reg[5]  ( .D(n718), .C(CLK_top), .QN(\position1/n365 ) );
  DF3 \position1/bi_reg[6]  ( .D(n717), .C(CLK_top), .QN(\position1/n364 ) );
  DF3 \position1/bi_reg[7]  ( .D(n716), .C(CLK_top), .QN(\position1/n363 ) );
  DF3 \position1/gi_reg[0]  ( .D(n731), .C(CLK_top), .Q(\position1/gi [0]), 
        .QN(\position1/n362 ) );
  DF3 \position1/gi_reg[1]  ( .D(n730), .C(CLK_top), .Q(\position1/gi [1]) );
  DF3 \position1/gi_reg[2]  ( .D(n729), .C(CLK_top), .Q(\position1/gi [2]), 
        .QN(\position1/n360 ) );
  DF3 \position1/gi_reg[3]  ( .D(n728), .C(CLK_top), .Q(\position1/gi [3]) );
  DF3 \position1/gi_reg[4]  ( .D(n727), .C(CLK_top), .Q(\position1/gi [4]), 
        .QN(\position1/n358 ) );
  DF3 \position1/gi_reg[5]  ( .D(n726), .C(CLK_top), .Q(\position1/gi [5]), 
        .QN(\position1/n357 ) );
  DF3 \position1/gi_reg[6]  ( .D(n725), .C(CLK_top), .Q(\position1/gi [6]), 
        .QN(\position1/n356 ) );
  DF3 \position1/gi_reg[7]  ( .D(n724), .C(CLK_top), .Q(\position1/gi [7]) );
  DF3 \position1/ri_reg[0]  ( .D(n739), .C(CLK_top), .QN(\position1/n353 ) );
  DF3 \position1/ri_reg[1]  ( .D(n738), .C(CLK_top), .QN(\position1/n352 ) );
  DF3 \position1/ri_reg[2]  ( .D(n737), .C(CLK_top), .QN(\position1/n351 ) );
  DF3 \position1/ri_reg[3]  ( .D(n736), .C(CLK_top), .QN(\position1/n350 ) );
  DF3 \position1/ri_reg[4]  ( .D(n735), .C(CLK_top), .QN(\position1/n349 ) );
  DF3 \position1/ri_reg[5]  ( .D(n734), .C(CLK_top), .QN(\position1/n348 ) );
  DF3 \position1/ri_reg[6]  ( .D(n733), .C(CLK_top), .QN(\position1/n347 ) );
  DF3 \position1/ri_reg[7]  ( .D(n732), .C(CLK_top), .QN(\position1/n346 ) );
  DFE1 \image_process1/r_out_reg[0]  ( .D(\image_process1/N8 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[0]) );
  DFE1 \image_process1/r_out_reg[1]  ( .D(\image_process1/N11 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[1]) );
  DFE1 \image_process1/r_out_reg[2]  ( .D(\image_process1/N14 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[2]) );
  DFE1 \image_process1/r_out_reg[3]  ( .D(\image_process1/N17 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[3]) );
  DFE1 \image_process1/r_out_reg[4]  ( .D(\image_process1/N20 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[4]) );
  DFE1 \image_process1/r_out_reg[5]  ( .D(\image_process1/N23 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[5]) );
  DFE1 \image_process1/r_out_reg[6]  ( .D(\image_process1/N26 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[6]) );
  DFE1 \image_process1/r_out_reg[7]  ( .D(\image_process1/N29 ), .E(reset_top), 
        .C(CLK_top), .Q(r_out_proc[7]) );
  DFE1 \image_process1/b_out_reg[0]  ( .D(\image_process1/N10 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[0]) );
  DFE1 \image_process1/b_out_reg[1]  ( .D(\image_process1/N13 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[1]) );
  DFE1 \image_process1/b_out_reg[2]  ( .D(\image_process1/N16 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[2]) );
  DFE1 \image_process1/b_out_reg[3]  ( .D(\image_process1/N19 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[3]) );
  DFE1 \image_process1/b_out_reg[4]  ( .D(\image_process1/N22 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[4]) );
  DFE1 \image_process1/b_out_reg[5]  ( .D(\image_process1/N25 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[5]) );
  DFE1 \image_process1/b_out_reg[6]  ( .D(\image_process1/N28 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[6]) );
  DFE1 \image_process1/b_out_reg[7]  ( .D(\image_process1/N31 ), .E(reset_top), 
        .C(CLK_top), .Q(b_out_proc[7]) );
  DFE1 \image_process1/g_out_reg[2]  ( .D(n767), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[2]) );
  DFE1 \image_process1/g_out_reg[6]  ( .D(n771), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[6]) );
  DFE1 \image_process1/g_out_reg[4]  ( .D(n769), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[4]) );
  DFE1 \image_process1/g_out_reg[5]  ( .D(n770), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[5]) );
  DFE1 \image_process1/g_out_reg[0]  ( .D(n773), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[0]) );
  DFE1 \image_process1/g_out_reg[1]  ( .D(n766), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[1]) );
  DFE1 \image_process1/g_out_reg[3]  ( .D(n768), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[3]) );
  DFE1 \image_process1/g_out_reg[7]  ( .D(n772), .E(reset_top), .C(CLK_top), 
        .Q(g_out_proc[7]) );
  XOR31 \position1/sub_226/U2_24  ( .A(\position1/y_sum [24]), .B(n44), .C(
        \position1/sub_226/carry [24]), .Q(\position1/N1962 ) );
  XOR31 \position1/sub_216/U2_24  ( .A(\position1/x_sum [24]), .B(n300), .C(
        \position1/sub_216/carry [24]), .Q(\position1/N1545 ) );
  XOR31 \position1/sub_226_I2/U2_24  ( .A(\position1/N1987 ), .B(n588), .C(
        \position1/sub_226_I2/carry [24]), .Q(\position1/N2014 ) );
  XOR31 \position1/sub_216_I2/U2_24  ( .A(\position1/N1570 ), .B(n589), .C(
        \position1/sub_216_I2/carry [24]), .Q(\position1/N1597 ) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_7  ( .A(n489), .B(
        cam_x[7]), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [7]), 
        .Q(\position1/dp_cluster_3/add_1_root_add_188_3/carry [8]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_3  ( .A(n497), .B(
        cam_x[3]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [3]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [4]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_5  ( .A(n493), .B(
        cam_x[5]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [5]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [6]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_5  ( .A(n493), .B(
        cam_x[5]), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [5]), 
        .Q(\position1/dp_cluster_3/add_1_root_add_188_3/carry [6]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_1  ( .A(n501), .B(
        cam_x[1]), .C(cam_x[0]), .Q(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [2]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_1  ( .A(n501), .B(
        cam_x[1]), .C(n503), .Q(
        \position1/dp_cluster_7/add_1_root_add_170_3/carry [2]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_3  ( .A(cam_x[3]), .B(
        n497), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [3]), .Q(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [4]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_2  ( .A(n499), .B(
        cam_x[2]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [2]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [3]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_2  ( .A(cam_x[2]), .B(
        n499), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [2]), .Q(
        \position1/dp_cluster_3/add_1_root_add_188_3/carry [3]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_6  ( .A(n491), .B(
        cam_x[6]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [6]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [7]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_6  ( .A(n491), .B(
        cam_x[6]), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [6]), 
        .Q(\position1/dp_cluster_3/add_1_root_add_188_3/carry [7]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_4  ( .A(n495), .B(
        cam_x[4]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [4]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [5]) );
  MAJ31 \position1/dp_cluster_3/add_1_root_add_188_3/U1_4  ( .A(n495), .B(
        cam_x[4]), .C(\position1/dp_cluster_3/add_1_root_add_188_3/carry [4]), 
        .Q(\position1/dp_cluster_3/add_1_root_add_188_3/carry [5]) );
  MAJ31 \position1/dp_cluster_7/add_1_root_add_170_3/U1_7  ( .A(n489), .B(
        cam_x[7]), .C(\position1/dp_cluster_7/add_1_root_add_170_3/carry [7]), 
        .Q(\position1/dp_cluster_7/add_1_root_add_170_3/carry [8]) );
  DFE1 \gensync1/comptY_reg[4]  ( .D(\gensync1/N60 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N169 ), .QN(n13) );
  DFE1 \gensync1/comptY_reg[3]  ( .D(\gensync1/N59 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N170 ), .QN(n11) );
  DFE1 \gensync1/comptY_reg[1]  ( .D(\gensync1/N57 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N172 ), .QN(n9) );
  DFE1 \gensync1/comptY_reg[2]  ( .D(\gensync1/N58 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N171 ), .QN(n8) );
  DFE1 \gensync1/comptY_reg[0]  ( .D(\gensync1/N56 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N173 ), .QN(n3) );
  DFE1 \gensync1/comptY_reg[5]  ( .D(\gensync1/N61 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N168 ) );
  DFE1 \gensync1/comptY_reg[6]  ( .D(\gensync1/N62 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N167 ) );
  DFE1 \gensync1/comptY_reg[7]  ( .D(\gensync1/N63 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N166 ) );
  DFE1 \gensync1/comptY_reg[8]  ( .D(\gensync1/N64 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/N165 ) );
  DFE1 \gensync1/comptY_reg[9]  ( .D(\gensync1/N65 ), .E(\gensync1/n107 ), .C(
        CLK_top), .Q(\gensync1/comptY[9] ) );
  XOR21 U2 ( .A(\position1/y_sum [9]), .B(\position1/r409/carry [9]), .Q(
        \position1/N364 ) );
  XOR21 U3 ( .A(\position1/x_sum [9]), .B(\position1/r406/carry [9]), .Q(
        \position1/N289 ) );
  NAND31 U4 ( .A(\position1/N267 ), .B(IMG_top), .C(\position1/n1389 ), .Q(
        \position1/n1062 ) );
  AOI221 U5 ( .A(n1125), .B(n547), .C(\position1/N1909 ), .D(n551), .Q(
        \position1/n1384 ) );
  AOI221 U6 ( .A(n906), .B(n581), .C(\position1/N2326 ), .D(n585), .Q(
        \position1/n1208 ) );
  NOR21 U7 ( .A(\gensync1/n102 ), .B(n113), .Q(\gensync1/N31 ) );
  NOR21 U8 ( .A(n507), .B(n112), .Q(\gensync1/N65 ) );
  XOR21 U9 ( .A(\position1/x_sum [20]), .B(\position1/r406/carry [20]), .Q(
        \position1/N300 ) );
  XOR21 U10 ( .A(\position1/x_sum [22]), .B(\position1/r406/carry [22]), .Q(
        \position1/N302 ) );
  XOR21 U11 ( .A(\position1/x_sum [21]), .B(\position1/r406/carry [21]), .Q(
        \position1/N301 ) );
  XOR21 U12 ( .A(\position1/x_sum [23]), .B(\position1/r406/carry [23]), .Q(
        \position1/N303 ) );
  XOR21 U13 ( .A(\position1/x_sum [14]), .B(\position1/r406/carry [14]), .Q(
        \position1/N294 ) );
  XOR21 U14 ( .A(\position1/x_sum [16]), .B(\position1/r406/carry [16]), .Q(
        \position1/N296 ) );
  XOR21 U15 ( .A(\position1/x_sum [18]), .B(\position1/r406/carry [18]), .Q(
        \position1/N298 ) );
  XOR21 U16 ( .A(\position1/y_sum [20]), .B(\position1/r409/carry [20]), .Q(
        \position1/N375 ) );
  XOR21 U17 ( .A(\position1/y_sum [22]), .B(\position1/r409/carry [22]), .Q(
        \position1/N377 ) );
  XOR21 U18 ( .A(\position1/x_sum [15]), .B(\position1/r406/carry [15]), .Q(
        \position1/N295 ) );
  XOR21 U19 ( .A(\position1/x_sum [17]), .B(\position1/r406/carry [17]), .Q(
        \position1/N297 ) );
  XOR21 U20 ( .A(\position1/y_sum [19]), .B(\position1/r409/carry [19]), .Q(
        \position1/N374 ) );
  XOR21 U21 ( .A(\position1/x_sum [19]), .B(\position1/r406/carry [19]), .Q(
        \position1/N299 ) );
  XOR21 U22 ( .A(\position1/y_sum [21]), .B(\position1/r409/carry [21]), .Q(
        \position1/N376 ) );
  XOR21 U23 ( .A(\position1/y_sum [23]), .B(\position1/r409/carry [23]), .Q(
        \position1/N378 ) );
  XOR21 U24 ( .A(\position1/x_sum [10]), .B(\position1/r406/carry [10]), .Q(
        \position1/N290 ) );
  XOR21 U25 ( .A(\position1/x_sum [12]), .B(\position1/r406/carry [12]), .Q(
        \position1/N292 ) );
  XOR21 U26 ( .A(\position1/y_sum [14]), .B(\position1/r409/carry [14]), .Q(
        \position1/N369 ) );
  XOR21 U27 ( .A(\position1/y_sum [16]), .B(\position1/r409/carry [16]), .Q(
        \position1/N371 ) );
  XOR21 U28 ( .A(\position1/y_sum [18]), .B(\position1/r409/carry [18]), .Q(
        \position1/N373 ) );
  XOR21 U29 ( .A(\position1/y_sum [13]), .B(\position1/r409/carry [13]), .Q(
        \position1/N368 ) );
  XOR21 U30 ( .A(\position1/x_sum [13]), .B(\position1/r406/carry [13]), .Q(
        \position1/N293 ) );
  XOR21 U31 ( .A(\position1/y_sum [15]), .B(\position1/r409/carry [15]), .Q(
        \position1/N370 ) );
  XOR21 U32 ( .A(\position1/y_sum [17]), .B(\position1/r409/carry [17]), .Q(
        \position1/N372 ) );
  XOR21 U33 ( .A(\position1/x_sum [11]), .B(\position1/r406/carry [11]), .Q(
        \position1/N291 ) );
  XOR21 U34 ( .A(\position1/y_sum [10]), .B(\position1/r409/carry [10]), .Q(
        \position1/N365 ) );
  XOR21 U35 ( .A(\position1/y_sum [12]), .B(\position1/r409/carry [12]), .Q(
        \position1/N367 ) );
  XOR21 U36 ( .A(\position1/y_sum [11]), .B(\position1/r409/carry [11]), .Q(
        \position1/N366 ) );
  OAI2111 U37 ( .A(n2), .B(n1710), .C(n1046), .D(\position1/n1333 ), .Q(
        \position1/N2040 ) );
  OAI2111 U38 ( .A(n2), .B(n2044), .C(n1265), .D(\position1/n1529 ), .Q(
        \position1/N1623 ) );
  INV3 U39 ( .A(n102), .Q(n1816) );
  INV3 U40 ( .A(n103), .Q(n1482) );
  INV3 U41 ( .A(n108), .Q(n2009) );
  INV3 U42 ( .A(n109), .Q(n1675) );
  INV3 U43 ( .A(n110), .Q(n2010) );
  INV3 U44 ( .A(n111), .Q(n1676) );
  BUF2 U45 ( .A(\position1/n1071 ), .Q(n476) );
  BUF2 U46 ( .A(n2126), .Q(\position1/dp_cluster_7/N314 ) );
  BUF2 U47 ( .A(\position1/N2457 ), .Q(n468) );
  BUF2 U48 ( .A(\position1/N2453 ), .Q(n471) );
  BUF2 U49 ( .A(\image_process1/n61 ), .Q(n488) );
  BUF2 U50 ( .A(\position1/N2449 ), .Q(n474) );
  BUF2 U51 ( .A(\position1/N2447 ), .Q(n475) );
  NOR40 U52 ( .A(n1388), .B(\image_process1/gi [5]), .C(\image_process1/gi [7]), .D(\image_process1/gi [6]), .Q(\image_process1/N59 ) );
  NAND22 U53 ( .A(\gensync1/N9 ), .B(n649), .Q(\gensync1/n102 ) );
  BUF2 U54 ( .A(\position1/N194 ), .Q(n484) );
  INV3 U55 ( .A(\position1/n1500 ), .Q(n1208) );
  INV3 U56 ( .A(\position1/n1304 ), .Q(n989) );
  INV3 U57 ( .A(\position1/n1517 ), .Q(n1226) );
  INV3 U58 ( .A(\position1/n1321 ), .Q(n1007) );
  INV3 U59 ( .A(\position1/n1515 ), .Q(n1224) );
  INV3 U60 ( .A(\position1/n1319 ), .Q(n1005) );
  INV3 U61 ( .A(\position1/n1513 ), .Q(n1222) );
  INV3 U62 ( .A(\position1/n1317 ), .Q(n1003) );
  INV3 U63 ( .A(\position1/n1511 ), .Q(n1220) );
  INV3 U64 ( .A(\position1/n1315 ), .Q(n1001) );
  INV3 U65 ( .A(\position1/n1509 ), .Q(n1218) );
  INV3 U66 ( .A(\position1/n1313 ), .Q(n999) );
  INV3 U67 ( .A(\position1/n1476 ), .Q(n1181) );
  INV3 U68 ( .A(\position1/n1280 ), .Q(n962) );
  INV3 U69 ( .A(\position1/n1519 ), .Q(n1229) );
  INV3 U70 ( .A(\position1/n1323 ), .Q(n1010) );
  INV3 U71 ( .A(\position1/n1443 ), .Q(n1143) );
  INV3 U72 ( .A(\position1/n1247 ), .Q(n924) );
  INV3 U73 ( .A(\position1/n1485 ), .Q(n1192) );
  INV3 U74 ( .A(\position1/n1289 ), .Q(n973) );
  INV3 U75 ( .A(\position1/n1469 ), .Q(n1174) );
  INV3 U76 ( .A(\position1/n1273 ), .Q(n955) );
  INV3 U77 ( .A(\position1/n1467 ), .Q(n1172) );
  INV3 U78 ( .A(\position1/n1271 ), .Q(n953) );
  INV3 U79 ( .A(\position1/n1465 ), .Q(n1170) );
  INV3 U80 ( .A(\position1/n1269 ), .Q(n951) );
  INV3 U81 ( .A(\position1/n1463 ), .Q(n1168) );
  INV3 U82 ( .A(\position1/n1267 ), .Q(n949) );
  INV3 U83 ( .A(\position1/n1461 ), .Q(n1166) );
  INV3 U84 ( .A(\position1/n1265 ), .Q(n947) );
  INV3 U85 ( .A(\position1/n1471 ), .Q(n1176) );
  INV3 U86 ( .A(\position1/n1275 ), .Q(n957) );
  INV3 U87 ( .A(\position1/n1495 ), .Q(n1203) );
  INV3 U88 ( .A(\position1/n1299 ), .Q(n984) );
  INV3 U89 ( .A(\position1/n1491 ), .Q(n1199) );
  INV3 U90 ( .A(\position1/n1295 ), .Q(n980) );
  INV3 U91 ( .A(\position1/n1489 ), .Q(n1197) );
  INV3 U92 ( .A(\position1/n1293 ), .Q(n978) );
  INV3 U93 ( .A(\position1/n1487 ), .Q(n1195) );
  INV3 U94 ( .A(\position1/n1291 ), .Q(n976) );
  INV3 U95 ( .A(\position1/n1445 ), .Q(n1146) );
  INV3 U96 ( .A(\position1/n1249 ), .Q(n927) );
  INV3 U97 ( .A(\position1/n1493 ), .Q(n1201) );
  INV3 U98 ( .A(\position1/n1297 ), .Q(n982) );
  NAND31 U99 ( .A(\position1/n1386 ), .B(\position1/n1384 ), .C(
        \position1/n1385 ), .Q(n102) );
  NAND31 U100 ( .A(\position1/n1210 ), .B(\position1/n1208 ), .C(
        \position1/n1209 ), .Q(n103) );
  NOR21 U101 ( .A(\position1/sub_216_I7/carry [23]), .B(n1160), .Q(n124) );
  NOR21 U102 ( .A(\position1/sub_226_I7/carry [23]), .B(n941), .Q(n140) );
  NOR21 U103 ( .A(\position1/sub_216_I6/carry [23]), .B(n1186), .Q(n120) );
  NOR21 U104 ( .A(\position1/sub_226_I6/carry [23]), .B(n967), .Q(n136) );
  INV3 U105 ( .A(n123), .Q(\position1/sub_216_I7/carry [23]) );
  NOR21 U106 ( .A(\position1/sub_216_I7/carry [22]), .B(n1161), .Q(n123) );
  INV3 U107 ( .A(n139), .Q(\position1/sub_226_I7/carry [23]) );
  NOR21 U108 ( .A(\position1/sub_226_I7/carry [22]), .B(n942), .Q(n139) );
  INV3 U109 ( .A(n127), .Q(\position1/sub_216_I8/carry [22]) );
  NOR21 U110 ( .A(\position1/sub_216_I8/carry [21]), .B(n1128), .Q(n127) );
  INV3 U111 ( .A(n143), .Q(\position1/sub_226_I8/carry [22]) );
  NOR21 U112 ( .A(\position1/sub_226_I8/carry [21]), .B(n909), .Q(n143) );
  INV3 U113 ( .A(n128), .Q(\position1/sub_216_I8/carry [23]) );
  NOR21 U114 ( .A(\position1/sub_216_I8/carry [22]), .B(n1127), .Q(n128) );
  INV3 U115 ( .A(n144), .Q(\position1/sub_226_I8/carry [23]) );
  NOR21 U116 ( .A(\position1/sub_226_I8/carry [22]), .B(n908), .Q(n144) );
  INV3 U117 ( .A(\position1/n1421 ), .Q(n1115) );
  INV3 U118 ( .A(\position1/n1225 ), .Q(n896) );
  INV3 U119 ( .A(\position1/N2397 ), .Q(n840) );
  INV3 U120 ( .A(\position1/N2399 ), .Q(n838) );
  INV3 U121 ( .A(\position1/N2376 ), .Q(n848) );
  AOI221 U122 ( .A(n533), .B(\position1/N1686 ), .C(n531), .D(
        \position1/N1659 ), .Q(\position1/n1519 ) );
  AOI221 U123 ( .A(n567), .B(\position1/N2103 ), .C(n565), .D(
        \position1/N2076 ), .Q(\position1/n1323 ) );
  AOI221 U124 ( .A(n545), .B(\position1/N1843 ), .C(n543), .D(n1173), .Q(
        \position1/n1443 ) );
  AOI221 U125 ( .A(n579), .B(\position1/N2260 ), .C(n577), .D(n954), .Q(
        \position1/n1247 ) );
  AOI221 U126 ( .A(n545), .B(\position1/N1841 ), .C(n543), .D(n1175), .Q(
        \position1/n1445 ) );
  AOI221 U127 ( .A(n579), .B(\position1/N2258 ), .C(n577), .D(n956), .Q(
        \position1/n1249 ) );
  AOI221 U128 ( .A(n538), .B(\position1/N1747 ), .C(n535), .D(n1219), .Q(
        \position1/n1485 ) );
  AOI221 U129 ( .A(n572), .B(\position1/N2164 ), .C(n569), .D(n1000), .Q(
        \position1/n1289 ) );
  AOI221 U130 ( .A(n1144), .B(n547), .C(\position1/N1894 ), .D(n549), .Q(
        \position1/n1419 ) );
  AOI221 U131 ( .A(n925), .B(n581), .C(\position1/N2311 ), .D(n583), .Q(
        \position1/n1223 ) );
  AOI221 U132 ( .A(n541), .B(\position1/N1790 ), .C(n539), .D(n1202), .Q(
        \position1/n1469 ) );
  AOI221 U133 ( .A(n575), .B(\position1/N2207 ), .C(n573), .D(n983), .Q(
        \position1/n1273 ) );
  AOI221 U134 ( .A(n541), .B(\position1/N1792 ), .C(n539), .D(n1200), .Q(
        \position1/n1467 ) );
  AOI221 U135 ( .A(n575), .B(\position1/N2209 ), .C(n573), .D(n981), .Q(
        \position1/n1271 ) );
  AOI221 U136 ( .A(n541), .B(\position1/N1794 ), .C(n539), .D(n1198), .Q(
        \position1/n1465 ) );
  AOI221 U137 ( .A(n575), .B(\position1/N2211 ), .C(n573), .D(n979), .Q(
        \position1/n1269 ) );
  AOI221 U138 ( .A(n542), .B(\position1/N1796 ), .C(n539), .D(n1196), .Q(
        \position1/n1463 ) );
  AOI221 U139 ( .A(n576), .B(\position1/N2213 ), .C(n573), .D(n977), .Q(
        \position1/n1267 ) );
  AOI221 U140 ( .A(n542), .B(\position1/N1798 ), .C(n539), .D(n1194), .Q(
        \position1/n1461 ) );
  AOI221 U141 ( .A(n576), .B(\position1/N2215 ), .C(n573), .D(n975), .Q(
        \position1/n1265 ) );
  AOI221 U142 ( .A(n541), .B(\position1/N1788 ), .C(n539), .D(n1204), .Q(
        \position1/n1471 ) );
  AOI221 U143 ( .A(n575), .B(\position1/N2205 ), .C(n573), .D(n985), .Q(
        \position1/n1275 ) );
  AOI221 U144 ( .A(n537), .B(\position1/N1737 ), .C(n535), .D(n1231), .Q(
        \position1/n1495 ) );
  AOI221 U145 ( .A(n571), .B(\position1/N2154 ), .C(n569), .D(n1012), .Q(
        \position1/n1299 ) );
  AOI221 U146 ( .A(n537), .B(\position1/N1741 ), .C(n535), .D(n1225), .Q(
        \position1/n1491 ) );
  AOI221 U147 ( .A(n571), .B(\position1/N2158 ), .C(n569), .D(n1006), .Q(
        \position1/n1295 ) );
  AOI221 U148 ( .A(n537), .B(\position1/N1743 ), .C(n535), .D(n1223), .Q(
        \position1/n1489 ) );
  AOI221 U149 ( .A(n571), .B(\position1/N2160 ), .C(n569), .D(n1004), .Q(
        \position1/n1293 ) );
  AOI221 U150 ( .A(n538), .B(\position1/N1745 ), .C(n535), .D(n1221), .Q(
        \position1/n1487 ) );
  AOI221 U151 ( .A(n572), .B(\position1/N2162 ), .C(n569), .D(n1002), .Q(
        \position1/n1291 ) );
  AOI221 U152 ( .A(n537), .B(\position1/N1739 ), .C(n535), .D(n1228), .Q(
        \position1/n1493 ) );
  AOI221 U153 ( .A(n571), .B(\position1/N2156 ), .C(n569), .D(n1009), .Q(
        \position1/n1297 ) );
  AOI221 U154 ( .A(n533), .B(\position1/N1688 ), .C(n531), .D(
        \position1/N1661 ), .Q(\position1/n1517 ) );
  AOI221 U155 ( .A(n567), .B(\position1/N2105 ), .C(n565), .D(
        \position1/N2078 ), .Q(\position1/n1321 ) );
  AOI221 U156 ( .A(n533), .B(\position1/N1690 ), .C(n531), .D(
        \position1/N1663 ), .Q(\position1/n1515 ) );
  AOI221 U157 ( .A(n567), .B(\position1/N2107 ), .C(n565), .D(
        \position1/N2080 ), .Q(\position1/n1319 ) );
  AOI221 U158 ( .A(n534), .B(\position1/N1692 ), .C(n531), .D(
        \position1/N1665 ), .Q(\position1/n1513 ) );
  AOI221 U159 ( .A(n568), .B(\position1/N2109 ), .C(n565), .D(
        \position1/N2082 ), .Q(\position1/n1317 ) );
  AOI221 U160 ( .A(n534), .B(\position1/N1694 ), .C(n531), .D(
        \position1/N1667 ), .Q(\position1/n1511 ) );
  AOI221 U161 ( .A(n568), .B(\position1/N2111 ), .C(n565), .D(
        \position1/N2084 ), .Q(\position1/n1315 ) );
  AOI221 U162 ( .A(n534), .B(\position1/N1696 ), .C(n531), .D(
        \position1/N1669 ), .Q(\position1/n1509 ) );
  AOI221 U163 ( .A(n568), .B(\position1/N2113 ), .C(n565), .D(
        \position1/N2086 ), .Q(\position1/n1313 ) );
  AOI221 U164 ( .A(n1142), .B(n547), .C(\position1/N1896 ), .D(n549), .Q(
        \position1/n1417 ) );
  AOI221 U165 ( .A(n923), .B(n581), .C(\position1/N2313 ), .D(n583), .Q(
        \position1/n1221 ) );
  AOI221 U166 ( .A(n1138), .B(n547), .C(\position1/N1898 ), .D(n550), .Q(
        \position1/n1415 ) );
  AOI221 U167 ( .A(n919), .B(n581), .C(\position1/N2315 ), .D(n584), .Q(
        \position1/n1219 ) );
  AOI221 U168 ( .A(n1135), .B(n547), .C(\position1/N1900 ), .D(n550), .Q(
        \position1/n1413 ) );
  AOI221 U169 ( .A(n916), .B(n581), .C(\position1/N2317 ), .D(n584), .Q(
        \position1/n1217 ) );
  AOI221 U170 ( .A(n536), .B(n1240), .C(n535), .D(n1240), .Q(\position1/n1500 ) );
  AOI221 U171 ( .A(n570), .B(n1021), .C(n569), .D(n1021), .Q(\position1/n1304 ) );
  AOI221 U172 ( .A(n1150), .B(n547), .C(\position1/N1890 ), .D(n549), .Q(
        \position1/n1423 ) );
  AOI221 U173 ( .A(n931), .B(n581), .C(\position1/N2307 ), .D(n583), .Q(
        \position1/n1227 ) );
  AOI221 U174 ( .A(n1147), .B(n547), .C(\position1/N1892 ), .D(n549), .Q(
        \position1/n1421 ) );
  AOI221 U175 ( .A(n928), .B(n581), .C(\position1/N2309 ), .D(n583), .Q(
        \position1/n1225 ) );
  AOI221 U176 ( .A(n540), .B(n1209), .C(n539), .D(n1209), .Q(\position1/n1476 ) );
  AOI221 U177 ( .A(n574), .B(n990), .C(n573), .D(n990), .Q(\position1/n1280 )
         );
  INV3 U178 ( .A(n548), .Q(n547) );
  INV3 U179 ( .A(n582), .Q(n581) );
  INV3 U180 ( .A(n544), .Q(n543) );
  INV3 U181 ( .A(n578), .Q(n577) );
  INV3 U182 ( .A(n540), .Q(n539) );
  INV3 U183 ( .A(n574), .Q(n573) );
  INV3 U184 ( .A(n532), .Q(n531) );
  INV3 U185 ( .A(n566), .Q(n565) );
  INV3 U186 ( .A(n536), .Q(n535) );
  INV3 U187 ( .A(n570), .Q(n569) );
  AOI221 U188 ( .A(n1126), .B(n547), .C(\position1/N1908 ), .D(n551), .Q(
        \position1/n1385 ) );
  XNR21 U189 ( .A(n1126), .B(\position1/sub_216_I8/carry [23]), .Q(
        \position1/N1908 ) );
  XOR21 U190 ( .A(n129), .B(n1125), .Q(\position1/N1909 ) );
  NOR21 U191 ( .A(\position1/sub_216_I8/carry [23]), .B(n1126), .Q(n129) );
  AOI221 U192 ( .A(n1127), .B(n547), .C(\position1/N1907 ), .D(n551), .Q(
        \position1/n1386 ) );
  XNR21 U193 ( .A(n1127), .B(\position1/sub_216_I8/carry [22]), .Q(
        \position1/N1907 ) );
  AOI221 U194 ( .A(n1128), .B(n547), .C(\position1/N1906 ), .D(n550), .Q(
        \position1/n1387 ) );
  XNR21 U195 ( .A(n1128), .B(\position1/sub_216_I8/carry [21]), .Q(
        \position1/N1906 ) );
  AOI221 U196 ( .A(n907), .B(n581), .C(\position1/N2325 ), .D(n585), .Q(
        \position1/n1209 ) );
  XNR21 U197 ( .A(n907), .B(\position1/sub_226_I8/carry [23]), .Q(
        \position1/N2325 ) );
  XOR21 U198 ( .A(n145), .B(n906), .Q(\position1/N2326 ) );
  NOR21 U199 ( .A(\position1/sub_226_I8/carry [23]), .B(n907), .Q(n145) );
  AOI221 U200 ( .A(n908), .B(n581), .C(\position1/N2324 ), .D(n585), .Q(
        \position1/n1210 ) );
  XNR21 U201 ( .A(n908), .B(\position1/sub_226_I8/carry [22]), .Q(
        \position1/N2324 ) );
  AOI221 U202 ( .A(n909), .B(n581), .C(\position1/N2323 ), .D(n584), .Q(
        \position1/n1211 ) );
  XNR21 U203 ( .A(n909), .B(\position1/sub_226_I8/carry [21]), .Q(
        \position1/N2323 ) );
  INV3 U204 ( .A(\position1/n1524 ), .Q(n1239) );
  INV3 U205 ( .A(\position1/n1328 ), .Q(n1020) );
  INV3 U206 ( .A(\position1/n1447 ), .Q(n1149) );
  AOI221 U207 ( .A(n545), .B(\position1/N1839 ), .C(n543), .D(n1177), .Q(
        \position1/n1447 ) );
  INV3 U208 ( .A(\position1/n1251 ), .Q(n930) );
  AOI221 U209 ( .A(n579), .B(\position1/N2256 ), .C(n577), .D(n958), .Q(
        \position1/n1251 ) );
  INV3 U210 ( .A(\position1/n1441 ), .Q(n1140) );
  AOI221 U211 ( .A(n545), .B(\position1/N1845 ), .C(n543), .D(n1171), .Q(
        \position1/n1441 ) );
  INV3 U212 ( .A(\position1/n1245 ), .Q(n921) );
  AOI221 U213 ( .A(n579), .B(\position1/N2262 ), .C(n577), .D(n952), .Q(
        \position1/n1245 ) );
  INV3 U214 ( .A(\position1/n1439 ), .Q(n1137) );
  AOI221 U215 ( .A(n545), .B(\position1/N1847 ), .C(n543), .D(n1169), .Q(
        \position1/n1439 ) );
  INV3 U216 ( .A(\position1/n1243 ), .Q(n918) );
  AOI221 U217 ( .A(n579), .B(\position1/N2264 ), .C(n577), .D(n950), .Q(
        \position1/n1243 ) );
  INV3 U218 ( .A(\position1/n1437 ), .Q(n1134) );
  AOI221 U219 ( .A(n546), .B(\position1/N1849 ), .C(n543), .D(n1167), .Q(
        \position1/n1437 ) );
  INV3 U220 ( .A(\position1/n1241 ), .Q(n915) );
  AOI221 U221 ( .A(n580), .B(\position1/N2266 ), .C(n577), .D(n948), .Q(
        \position1/n1241 ) );
  INV3 U222 ( .A(n528), .Q(n526) );
  INV3 U223 ( .A(n562), .Q(n560) );
  INV3 U224 ( .A(\position1/n1516 ), .Q(n1225) );
  INV3 U225 ( .A(\position1/n1320 ), .Q(n1006) );
  INV3 U226 ( .A(\position1/n1514 ), .Q(n1223) );
  INV3 U227 ( .A(\position1/n1318 ), .Q(n1004) );
  INV3 U228 ( .A(\position1/n1512 ), .Q(n1221) );
  INV3 U229 ( .A(\position1/n1316 ), .Q(n1002) );
  INV3 U230 ( .A(\position1/n1510 ), .Q(n1219) );
  INV3 U231 ( .A(\position1/n1314 ), .Q(n1000) );
  INV3 U232 ( .A(\position1/n1508 ), .Q(n1217) );
  INV3 U233 ( .A(\position1/n1312 ), .Q(n998) );
  INV3 U234 ( .A(\position1/n1456 ), .Q(n1161) );
  AOI221 U235 ( .A(n542), .B(\position1/N1803 ), .C(n539), .D(n1187), .Q(
        \position1/n1456 ) );
  XNR21 U236 ( .A(n1187), .B(\position1/sub_216_I6/carry [22]), .Q(
        \position1/N1803 ) );
  INV3 U237 ( .A(\position1/n1260 ), .Q(n942) );
  AOI221 U238 ( .A(n576), .B(\position1/N2220 ), .C(n573), .D(n968), .Q(
        \position1/n1260 ) );
  XNR21 U239 ( .A(n968), .B(\position1/sub_226_I6/carry [22]), .Q(
        \position1/N2220 ) );
  INV3 U240 ( .A(\position1/n1455 ), .Q(n1160) );
  AOI221 U241 ( .A(n542), .B(\position1/N1804 ), .C(n539), .D(n1186), .Q(
        \position1/n1455 ) );
  XNR21 U242 ( .A(n1186), .B(\position1/sub_216_I6/carry [23]), .Q(
        \position1/N1804 ) );
  INV3 U243 ( .A(\position1/n1259 ), .Q(n941) );
  AOI221 U244 ( .A(n576), .B(\position1/N2221 ), .C(n573), .D(n967), .Q(
        \position1/n1259 ) );
  XNR21 U245 ( .A(n967), .B(\position1/sub_226_I6/carry [23]), .Q(
        \position1/N2221 ) );
  INV3 U246 ( .A(\position1/n1460 ), .Q(n1165) );
  INV3 U247 ( .A(\position1/n1264 ), .Q(n946) );
  INV3 U248 ( .A(\position1/n1494 ), .Q(n1202) );
  INV3 U249 ( .A(\position1/n1298 ), .Q(n983) );
  INV3 U250 ( .A(\position1/n1492 ), .Q(n1200) );
  INV3 U251 ( .A(\position1/n1296 ), .Q(n981) );
  INV3 U252 ( .A(\position1/n1490 ), .Q(n1198) );
  INV3 U253 ( .A(\position1/n1294 ), .Q(n979) );
  INV3 U254 ( .A(\position1/n1488 ), .Q(n1196) );
  INV3 U255 ( .A(\position1/n1292 ), .Q(n977) );
  INV3 U256 ( .A(\position1/n1486 ), .Q(n1194) );
  INV3 U257 ( .A(\position1/n1290 ), .Q(n975) );
  INV3 U258 ( .A(\position1/n1498 ), .Q(n1206) );
  INV3 U259 ( .A(\position1/n1302 ), .Q(n987) );
  INV3 U260 ( .A(\position1/n1496 ), .Q(n1204) );
  INV3 U261 ( .A(\position1/n1300 ), .Q(n985) );
  INV3 U262 ( .A(\position1/n1432 ), .Q(n1128) );
  AOI221 U263 ( .A(n546), .B(\position1/N1854 ), .C(n543), .D(n1162), .Q(
        \position1/n1432 ) );
  XNR21 U264 ( .A(n1162), .B(\position1/sub_216_I7/carry [21]), .Q(
        \position1/N1854 ) );
  INV3 U265 ( .A(\position1/n1431 ), .Q(n1127) );
  AOI221 U266 ( .A(n546), .B(\position1/N1855 ), .C(n543), .D(n1161), .Q(
        \position1/n1431 ) );
  XNR21 U267 ( .A(n1161), .B(\position1/sub_216_I7/carry [22]), .Q(
        \position1/N1855 ) );
  INV3 U268 ( .A(\position1/n1236 ), .Q(n909) );
  AOI221 U269 ( .A(n580), .B(\position1/N2271 ), .C(n577), .D(n943), .Q(
        \position1/n1236 ) );
  XNR21 U270 ( .A(n943), .B(\position1/sub_226_I7/carry [21]), .Q(
        \position1/N2271 ) );
  INV3 U271 ( .A(\position1/n1235 ), .Q(n908) );
  AOI221 U272 ( .A(n580), .B(\position1/N2272 ), .C(n577), .D(n942), .Q(
        \position1/n1235 ) );
  XNR21 U273 ( .A(n942), .B(\position1/sub_226_I7/carry [22]), .Q(
        \position1/N2272 ) );
  INV3 U274 ( .A(\position1/n1430 ), .Q(n1126) );
  AOI221 U275 ( .A(n546), .B(\position1/N1856 ), .C(n543), .D(n1160), .Q(
        \position1/n1430 ) );
  XNR21 U276 ( .A(n1160), .B(\position1/sub_216_I7/carry [23]), .Q(
        \position1/N1856 ) );
  INV3 U277 ( .A(\position1/n1234 ), .Q(n907) );
  AOI221 U278 ( .A(n580), .B(\position1/N2273 ), .C(n577), .D(n941), .Q(
        \position1/n1234 ) );
  XNR21 U279 ( .A(n941), .B(\position1/sub_226_I7/carry [23]), .Q(
        \position1/N2273 ) );
  INV3 U280 ( .A(\position1/n1459 ), .Q(n1164) );
  INV3 U281 ( .A(\position1/n1263 ), .Q(n945) );
  INV3 U282 ( .A(\position1/n1520 ), .Q(n1231) );
  INV3 U283 ( .A(\position1/n1324 ), .Q(n1012) );
  INV3 U284 ( .A(\position1/n1473 ), .Q(n1178) );
  INV3 U285 ( .A(\position1/n1277 ), .Q(n959) );
  INV3 U286 ( .A(\position1/n1480 ), .Q(n1186) );
  AOI221 U287 ( .A(n538), .B(\position1/N1752 ), .C(n535), .D(n1214), .Q(
        \position1/n1480 ) );
  XNR21 U288 ( .A(n1214), .B(\position1/sub_216_I5/carry [23]), .Q(
        \position1/N1752 ) );
  INV3 U289 ( .A(\position1/n1284 ), .Q(n967) );
  AOI221 U290 ( .A(n572), .B(\position1/N2169 ), .C(n569), .D(n995), .Q(
        \position1/n1284 ) );
  XNR21 U291 ( .A(n995), .B(\position1/sub_226_I5/carry [23]), .Q(
        \position1/N2169 ) );
  INV3 U292 ( .A(\position1/n1522 ), .Q(n1235) );
  INV3 U293 ( .A(\position1/n1326 ), .Q(n1016) );
  INV3 U294 ( .A(\position1/n1435 ), .Q(n1132) );
  INV3 U295 ( .A(\position1/n1239 ), .Q(n913) );
  INV3 U296 ( .A(\position1/n1497 ), .Q(n1205) );
  INV3 U297 ( .A(\position1/n1301 ), .Q(n986) );
  INV3 U298 ( .A(n528), .Q(n527) );
  INV3 U299 ( .A(n562), .Q(n561) );
  INV3 U300 ( .A(\position1/n1452 ), .Q(n1157) );
  AOI221 U301 ( .A(n544), .B(n1182), .C(n543), .D(n1182), .Q(\position1/n1452 ) );
  INV3 U302 ( .A(\position1/n1256 ), .Q(n938) );
  AOI221 U303 ( .A(n578), .B(n963), .C(n577), .D(n963), .Q(\position1/n1256 )
         );
  INV3 U304 ( .A(\position1/n1436 ), .Q(n1133) );
  INV3 U305 ( .A(\position1/n1240 ), .Q(n914) );
  INV3 U306 ( .A(\position1/n1474 ), .Q(n1179) );
  INV3 U307 ( .A(\position1/n1278 ), .Q(n960) );
  INV3 U308 ( .A(\position1/n1472 ), .Q(n1177) );
  INV3 U309 ( .A(\position1/n1276 ), .Q(n958) );
  INV3 U310 ( .A(\position1/n1470 ), .Q(n1175) );
  INV3 U311 ( .A(\position1/n1274 ), .Q(n956) );
  INV3 U312 ( .A(\position1/n1466 ), .Q(n1171) );
  INV3 U313 ( .A(\position1/n1270 ), .Q(n952) );
  INV3 U314 ( .A(\position1/n1464 ), .Q(n1169) );
  INV3 U315 ( .A(\position1/n1268 ), .Q(n950) );
  INV3 U316 ( .A(\position1/n1462 ), .Q(n1167) );
  INV3 U317 ( .A(\position1/n1266 ), .Q(n948) );
  INV3 U318 ( .A(\position1/n1468 ), .Q(n1173) );
  INV3 U319 ( .A(\position1/n1272 ), .Q(n954) );
  INV3 U320 ( .A(\position1/n1507 ), .Q(n1216) );
  INV3 U321 ( .A(\position1/n1311 ), .Q(n997) );
  INV3 U322 ( .A(\position1/n1450 ), .Q(n1153) );
  INV3 U323 ( .A(\position1/n1254 ), .Q(n934) );
  INV3 U324 ( .A(\position1/n1448 ), .Q(n1150) );
  INV3 U325 ( .A(\position1/n1252 ), .Q(n931) );
  INV3 U326 ( .A(\position1/n1446 ), .Q(n1147) );
  INV3 U327 ( .A(\position1/n1250 ), .Q(n928) );
  INV3 U328 ( .A(\position1/n1440 ), .Q(n1138) );
  INV3 U329 ( .A(\position1/n1244 ), .Q(n919) );
  INV3 U330 ( .A(\position1/n1438 ), .Q(n1135) );
  INV3 U331 ( .A(\position1/n1242 ), .Q(n916) );
  INV3 U332 ( .A(\position1/n1454 ), .Q(n1159) );
  AOI221 U333 ( .A(n542), .B(\position1/N1805 ), .C(n539), .D(n1185), .Q(
        \position1/n1454 ) );
  XNR21 U334 ( .A(\position1/sub_216_I6/carry [24]), .B(n1185), .Q(
        \position1/N1805 ) );
  INV3 U335 ( .A(n120), .Q(\position1/sub_216_I6/carry [24]) );
  INV3 U336 ( .A(\position1/n1258 ), .Q(n940) );
  AOI221 U337 ( .A(n576), .B(\position1/N2222 ), .C(n573), .D(n966), .Q(
        \position1/n1258 ) );
  XNR21 U338 ( .A(\position1/sub_226_I6/carry [24]), .B(n966), .Q(
        \position1/N2222 ) );
  INV3 U339 ( .A(n136), .Q(\position1/sub_226_I6/carry [24]) );
  INV3 U340 ( .A(\position1/n1429 ), .Q(n1125) );
  AOI221 U341 ( .A(n546), .B(\position1/N1857 ), .C(n543), .D(n1159), .Q(
        \position1/n1429 ) );
  XNR21 U342 ( .A(\position1/sub_216_I7/carry [24]), .B(n1159), .Q(
        \position1/N1857 ) );
  INV3 U343 ( .A(n124), .Q(\position1/sub_216_I7/carry [24]) );
  INV3 U344 ( .A(\position1/n1233 ), .Q(n906) );
  AOI221 U345 ( .A(n580), .B(\position1/N2274 ), .C(n577), .D(n940), .Q(
        \position1/n1233 ) );
  XNR21 U346 ( .A(\position1/sub_226_I7/carry [24]), .B(n940), .Q(
        \position1/N2274 ) );
  INV3 U347 ( .A(n140), .Q(\position1/sub_226_I7/carry [24]) );
  INV3 U348 ( .A(\position1/n1479 ), .Q(n1185) );
  AOI221 U349 ( .A(n538), .B(\position1/N1753 ), .C(n535), .D(n1213), .Q(
        \position1/n1479 ) );
  XNR21 U350 ( .A(\position1/sub_216_I5/carry [24]), .B(n1213), .Q(
        \position1/N1753 ) );
  INV3 U351 ( .A(n117), .Q(\position1/sub_216_I5/carry [24]) );
  INV3 U352 ( .A(\position1/n1283 ), .Q(n966) );
  AOI221 U353 ( .A(n572), .B(\position1/N2170 ), .C(n569), .D(n994), .Q(
        \position1/n1283 ) );
  XNR21 U354 ( .A(\position1/sub_226_I5/carry [24]), .B(n994), .Q(
        \position1/N2170 ) );
  INV3 U355 ( .A(n133), .Q(\position1/sub_226_I5/carry [24]) );
  INV3 U356 ( .A(\position1/n1453 ), .Q(n1158) );
  AOI221 U357 ( .A(n544), .B(n1183), .C(n543), .D(n1183), .Q(\position1/n1453 ) );
  INV3 U358 ( .A(\position1/n1257 ), .Q(n939) );
  AOI221 U359 ( .A(n578), .B(n964), .C(n577), .D(n964), .Q(\position1/n1257 )
         );
  INV3 U360 ( .A(\position1/n1502 ), .Q(n1210) );
  AOI221 U361 ( .A(n536), .B(n1242), .C(n535), .D(n1242), .Q(\position1/n1502 ) );
  INV3 U362 ( .A(\position1/n1501 ), .Q(n1209) );
  AOI221 U363 ( .A(n536), .B(n1241), .C(n535), .D(n1241), .Q(\position1/n1501 ) );
  INV3 U364 ( .A(\position1/n1503 ), .Q(n1211) );
  AOI221 U365 ( .A(n536), .B(n1243), .C(n535), .D(n1243), .Q(\position1/n1503 ) );
  INV3 U366 ( .A(\position1/n1306 ), .Q(n991) );
  AOI221 U367 ( .A(n570), .B(n1023), .C(n569), .D(n1023), .Q(\position1/n1306 ) );
  INV3 U368 ( .A(\position1/n1305 ), .Q(n990) );
  AOI221 U369 ( .A(n570), .B(n1022), .C(n569), .D(n1022), .Q(\position1/n1305 ) );
  INV3 U370 ( .A(\position1/n1307 ), .Q(n992) );
  AOI221 U371 ( .A(n570), .B(n1024), .C(n569), .D(n1024), .Q(\position1/n1307 ) );
  INV3 U372 ( .A(\position1/n1478 ), .Q(n1183) );
  AOI221 U373 ( .A(n540), .B(n1211), .C(n539), .D(n1211), .Q(\position1/n1478 ) );
  INV3 U374 ( .A(\position1/n1477 ), .Q(n1182) );
  AOI221 U375 ( .A(n540), .B(n1210), .C(n539), .D(n1210), .Q(\position1/n1477 ) );
  INV3 U376 ( .A(\position1/n1282 ), .Q(n964) );
  AOI221 U377 ( .A(n574), .B(n992), .C(n573), .D(n992), .Q(\position1/n1282 )
         );
  INV3 U378 ( .A(\position1/n1281 ), .Q(n963) );
  AOI221 U379 ( .A(n574), .B(n991), .C(n573), .D(n991), .Q(\position1/n1281 )
         );
  NOR21 U380 ( .A(\position1/sub_216_I5/carry [23]), .B(n1214), .Q(n117) );
  NOR21 U381 ( .A(\position1/sub_226_I5/carry [23]), .B(n995), .Q(n133) );
  XNR21 U382 ( .A(n1129), .B(\position1/sub_216_I8/carry [20]), .Q(
        \position1/N1905 ) );
  XNR21 U383 ( .A(n910), .B(\position1/sub_226_I8/carry [20]), .Q(
        \position1/N2322 ) );
  BUF2 U384 ( .A(n530), .Q(n529) );
  BUF2 U385 ( .A(n564), .Q(n563) );
  INV3 U386 ( .A(n119), .Q(\position1/sub_216_I6/carry [23]) );
  NOR21 U387 ( .A(\position1/sub_216_I6/carry [22]), .B(n1187), .Q(n119) );
  INV3 U388 ( .A(n135), .Q(\position1/sub_226_I6/carry [23]) );
  NOR21 U389 ( .A(\position1/sub_226_I6/carry [22]), .B(n968), .Q(n135) );
  INV3 U390 ( .A(n122), .Q(\position1/sub_216_I7/carry [22]) );
  NOR21 U391 ( .A(\position1/sub_216_I7/carry [21]), .B(n1162), .Q(n122) );
  INV3 U392 ( .A(n126), .Q(\position1/sub_216_I8/carry [21]) );
  NOR21 U393 ( .A(\position1/sub_216_I8/carry [20]), .B(n1129), .Q(n126) );
  INV3 U394 ( .A(n138), .Q(\position1/sub_226_I7/carry [22]) );
  NOR21 U395 ( .A(\position1/sub_226_I7/carry [21]), .B(n943), .Q(n138) );
  INV3 U396 ( .A(n142), .Q(\position1/sub_226_I8/carry [21]) );
  NOR21 U397 ( .A(\position1/sub_226_I8/carry [20]), .B(n910), .Q(n142) );
  INV3 U398 ( .A(\position1/n1416 ), .Q(n1109) );
  INV3 U399 ( .A(\position1/n1220 ), .Q(n890) );
  INV3 U400 ( .A(\position1/n1414 ), .Q(n1107) );
  INV3 U401 ( .A(\position1/n1218 ), .Q(n888) );
  INV3 U402 ( .A(\position1/n1426 ), .Q(n1120) );
  INV3 U403 ( .A(\position1/n1230 ), .Q(n901) );
  INV3 U404 ( .A(\position1/n1424 ), .Q(n1118) );
  INV3 U405 ( .A(\position1/n1228 ), .Q(n899) );
  INV3 U406 ( .A(\position1/n1422 ), .Q(n1116) );
  INV3 U407 ( .A(\position1/n1226 ), .Q(n897) );
  NOR21 U408 ( .A(n1101), .B(n1102), .Q(n1817) );
  INV3 U409 ( .A(\position1/n1388 ), .Q(n1102) );
  INV3 U410 ( .A(\position1/n1387 ), .Q(n1101) );
  AOI221 U411 ( .A(n1129), .B(n547), .C(\position1/N1905 ), .D(n550), .Q(
        \position1/n1388 ) );
  NOR21 U412 ( .A(n882), .B(n883), .Q(n1483) );
  INV3 U413 ( .A(\position1/n1212 ), .Q(n883) );
  INV3 U414 ( .A(\position1/n1211 ), .Q(n882) );
  AOI221 U415 ( .A(n910), .B(n581), .C(\position1/N2322 ), .D(n584), .Q(
        \position1/n1212 ) );
  INV3 U416 ( .A(\position1/n1428 ), .Q(n1122) );
  AOI221 U417 ( .A(n1158), .B(n547), .C(n1158), .D(n548), .Q(\position1/n1428 ) );
  INV3 U418 ( .A(\position1/n1232 ), .Q(n903) );
  AOI221 U419 ( .A(n939), .B(n581), .C(n939), .D(n582), .Q(\position1/n1232 )
         );
  XOR21 U420 ( .A(n495), .B(\position1/add_250/carry[4] ), .Q(
        \position1/N2397 ) );
  XOR21 U421 ( .A(n491), .B(\position1/add_250/carry[6] ), .Q(
        \position1/N2399 ) );
  XNR21 U422 ( .A(n495), .B(\position1/sub_250/carry[4] ), .Q(
        \position1/N2376 ) );
  XNR21 U423 ( .A(n491), .B(\position1/sub_250/carry[6] ), .Q(
        \position1/N2378 ) );
  BUF2 U424 ( .A(\position1/n856 ), .Q(n637) );
  BUF2 U425 ( .A(\position1/n856 ), .Q(n636) );
  BUF2 U426 ( .A(\position1/n856 ), .Q(n635) );
  NAND22 U427 ( .A(n741), .B(n782), .Q(\position1/n1057 ) );
  BUF2 U428 ( .A(n740), .Q(n511) );
  BUF2 U429 ( .A(n740), .Q(n512) );
  INV3 U430 ( .A(n148), .Q(\position1/sub_250/carry[5] ) );
  NOR21 U431 ( .A(\position1/sub_250/carry[4] ), .B(n495), .Q(n148) );
  INV3 U432 ( .A(n150), .Q(\position1/sub_250/carry[7] ) );
  NOR21 U433 ( .A(\position1/sub_250/carry[6] ), .B(n491), .Q(n150) );
  INV3 U434 ( .A(\position1/N2409 ), .Q(n793) );
  INV3 U435 ( .A(\position1/N2398 ), .Q(n839) );
  INV3 U436 ( .A(\position1/N2400 ), .Q(n837) );
  INV3 U437 ( .A(\position1/N2377 ), .Q(n847) );
  INV3 U438 ( .A(\position1/N2379 ), .Q(n845) );
  NOR21 U439 ( .A(n311), .B(n312), .Q(\position1/add_250/carry[7] ) );
  INV3 U440 ( .A(n491), .Q(n312) );
  INV3 U441 ( .A(\position1/add_250/carry[6] ), .Q(n311) );
  NOR21 U442 ( .A(n307), .B(n308), .Q(\position1/add_250/carry[5] ) );
  INV3 U443 ( .A(n495), .Q(n308) );
  INV3 U444 ( .A(\position1/add_250/carry[4] ), .Q(n307) );
  BUF2 U445 ( .A(\position1/n859 ), .Q(n645) );
  BUF2 U446 ( .A(\position1/n859 ), .Q(n646) );
  BUF2 U447 ( .A(\position1/n859 ), .Q(n647) );
  BUF2 U448 ( .A(\position1/n856 ), .Q(n638) );
  INV3 U449 ( .A(\image_process1/n97 ), .Q(n776) );
  INV3 U450 ( .A(\position1/N1634 ), .Q(n1292) );
  INV3 U451 ( .A(\position1/N2051 ), .Q(n1073) );
  INV3 U452 ( .A(\position1/N1636 ), .Q(n1287) );
  INV3 U453 ( .A(\position1/N2053 ), .Q(n1068) );
  INV3 U454 ( .A(\position1/N1638 ), .Q(n1283) );
  INV3 U455 ( .A(\position1/N2055 ), .Q(n1064) );
  INV3 U456 ( .A(\position1/N1640 ), .Q(n1279) );
  INV3 U457 ( .A(\position1/N2057 ), .Q(n1060) );
  INV3 U458 ( .A(\position1/N1642 ), .Q(n1275) );
  INV3 U459 ( .A(\position1/N2059 ), .Q(n1056) );
  INV3 U460 ( .A(\position1/N1644 ), .Q(n1271) );
  INV3 U461 ( .A(\position1/N2061 ), .Q(n1052) );
  INV3 U462 ( .A(\position1/N1646 ), .Q(n1248) );
  INV3 U463 ( .A(\position1/N2063 ), .Q(n1029) );
  INV3 U464 ( .A(\position1/N1648 ), .Q(n1245) );
  INV3 U465 ( .A(\position1/N2065 ), .Q(n1026) );
  AOI221 U466 ( .A(n542), .B(\position1/N1799 ), .C(n539), .D(n1192), .Q(
        \position1/n1460 ) );
  AOI221 U467 ( .A(n576), .B(\position1/N2216 ), .C(n573), .D(n973), .Q(
        \position1/n1264 ) );
  AOI221 U468 ( .A(n546), .B(\position1/N1851 ), .C(n543), .D(n1165), .Q(
        \position1/n1435 ) );
  AOI221 U469 ( .A(n580), .B(\position1/N2268 ), .C(n577), .D(n946), .Q(
        \position1/n1239 ) );
  AOI221 U470 ( .A(n542), .B(\position1/N1800 ), .C(n539), .D(n1191), .Q(
        \position1/n1459 ) );
  AOI221 U471 ( .A(n576), .B(\position1/N2217 ), .C(n573), .D(n972), .Q(
        \position1/n1263 ) );
  AOI221 U472 ( .A(n533), .B(\position1/N1685 ), .C(n531), .D(
        \position1/N1658 ), .Q(\position1/n1520 ) );
  AOI221 U473 ( .A(n567), .B(\position1/N2102 ), .C(n565), .D(
        \position1/N2075 ), .Q(\position1/n1324 ) );
  AOI221 U474 ( .A(n533), .B(\position1/N1683 ), .C(n531), .D(
        \position1/N1656 ), .Q(\position1/n1522 ) );
  AOI221 U475 ( .A(n567), .B(\position1/N2100 ), .C(n565), .D(
        \position1/N2073 ), .Q(\position1/n1326 ) );
  AOI221 U476 ( .A(n546), .B(\position1/N1850 ), .C(n543), .D(n1166), .Q(
        \position1/n1436 ) );
  AOI221 U477 ( .A(n580), .B(\position1/N2267 ), .C(n577), .D(n947), .Q(
        \position1/n1240 ) );
  AOI221 U478 ( .A(n533), .B(\position1/N1654 ), .C(n531), .D(
        \position1/N1654 ), .Q(\position1/n1524 ) );
  AOI221 U479 ( .A(n567), .B(\position1/N2071 ), .C(n565), .D(
        \position1/N2071 ), .Q(\position1/n1328 ) );
  AOI221 U480 ( .A(n541), .B(\position1/N1786 ), .C(n539), .D(n1206), .Q(
        \position1/n1473 ) );
  AOI221 U481 ( .A(n575), .B(\position1/N2203 ), .C(n573), .D(n987), .Q(
        \position1/n1277 ) );
  AOI221 U482 ( .A(n537), .B(\position1/N1735 ), .C(n535), .D(n1235), .Q(
        \position1/n1497 ) );
  AOI221 U483 ( .A(n571), .B(\position1/N2152 ), .C(n569), .D(n1016), .Q(
        \position1/n1301 ) );
  AOI221 U484 ( .A(n1140), .B(n547), .C(\position1/N1897 ), .D(n549), .Q(
        \position1/n1416 ) );
  AOI221 U485 ( .A(n921), .B(n581), .C(\position1/N2314 ), .D(n583), .Q(
        \position1/n1220 ) );
  AOI221 U486 ( .A(n1137), .B(n547), .C(\position1/N1899 ), .D(n550), .Q(
        \position1/n1414 ) );
  AOI221 U487 ( .A(n918), .B(n581), .C(\position1/N2316 ), .D(n584), .Q(
        \position1/n1218 ) );
  AOI221 U488 ( .A(n1134), .B(n547), .C(\position1/N1901 ), .D(n550), .Q(
        \position1/n1412 ) );
  AOI221 U489 ( .A(n915), .B(n581), .C(\position1/N2318 ), .D(n584), .Q(
        \position1/n1216 ) );
  AOI221 U490 ( .A(n1155), .B(n547), .C(\position1/N1887 ), .D(n548), .Q(
        \position1/n1426 ) );
  AOI221 U491 ( .A(n936), .B(n581), .C(\position1/N2304 ), .D(n582), .Q(
        \position1/n1230 ) );
  AOI221 U492 ( .A(n1152), .B(n547), .C(\position1/N1889 ), .D(n549), .Q(
        \position1/n1424 ) );
  AOI221 U493 ( .A(n933), .B(n581), .C(\position1/N2306 ), .D(n583), .Q(
        \position1/n1228 ) );
  AOI221 U494 ( .A(n1149), .B(n547), .C(\position1/N1891 ), .D(n549), .Q(
        \position1/n1422 ) );
  AOI221 U495 ( .A(n930), .B(n581), .C(\position1/N2308 ), .D(n583), .Q(
        \position1/n1226 ) );
  AOI221 U496 ( .A(n534), .B(\position1/N1698 ), .C(n531), .D(
        \position1/N1671 ), .Q(\position1/n1507 ) );
  AOI221 U497 ( .A(n568), .B(\position1/N2115 ), .C(n565), .D(
        \position1/N2088 ), .Q(\position1/n1311 ) );
  AOI221 U498 ( .A(n533), .B(\position1/N1689 ), .C(n531), .D(
        \position1/N1662 ), .Q(\position1/n1516 ) );
  AOI221 U499 ( .A(n567), .B(\position1/N2106 ), .C(n565), .D(
        \position1/N2079 ), .Q(\position1/n1320 ) );
  AOI221 U500 ( .A(n533), .B(\position1/N1691 ), .C(n531), .D(
        \position1/N1664 ), .Q(\position1/n1514 ) );
  AOI221 U501 ( .A(n567), .B(\position1/N2108 ), .C(n565), .D(
        \position1/N2081 ), .Q(\position1/n1318 ) );
  AOI221 U502 ( .A(n534), .B(\position1/N1693 ), .C(n531), .D(
        \position1/N1666 ), .Q(\position1/n1512 ) );
  AOI221 U503 ( .A(n568), .B(\position1/N2110 ), .C(n565), .D(
        \position1/N2083 ), .Q(\position1/n1316 ) );
  AOI221 U504 ( .A(n534), .B(\position1/N1695 ), .C(n531), .D(
        \position1/N1668 ), .Q(\position1/n1510 ) );
  AOI221 U505 ( .A(n568), .B(\position1/N2112 ), .C(n565), .D(
        \position1/N2085 ), .Q(\position1/n1314 ) );
  AOI221 U506 ( .A(n534), .B(\position1/N1697 ), .C(n531), .D(
        \position1/N1670 ), .Q(\position1/n1508 ) );
  AOI221 U507 ( .A(n568), .B(\position1/N2114 ), .C(n565), .D(
        \position1/N2087 ), .Q(\position1/n1312 ) );
  AOI221 U508 ( .A(n541), .B(\position1/N1785 ), .C(n539), .D(n1207), .Q(
        \position1/n1474 ) );
  AOI221 U509 ( .A(n575), .B(\position1/N2202 ), .C(n573), .D(n988), .Q(
        \position1/n1278 ) );
  AOI221 U510 ( .A(n541), .B(\position1/N1787 ), .C(n539), .D(n1205), .Q(
        \position1/n1472 ) );
  AOI221 U511 ( .A(n575), .B(\position1/N2204 ), .C(n573), .D(n986), .Q(
        \position1/n1276 ) );
  AOI221 U512 ( .A(n541), .B(\position1/N1789 ), .C(n539), .D(n1203), .Q(
        \position1/n1470 ) );
  AOI221 U513 ( .A(n575), .B(\position1/N2206 ), .C(n573), .D(n984), .Q(
        \position1/n1274 ) );
  AOI221 U514 ( .A(n541), .B(\position1/N1793 ), .C(n539), .D(n1199), .Q(
        \position1/n1466 ) );
  AOI221 U515 ( .A(n575), .B(\position1/N2210 ), .C(n573), .D(n980), .Q(
        \position1/n1270 ) );
  AOI221 U516 ( .A(n541), .B(\position1/N1795 ), .C(n539), .D(n1197), .Q(
        \position1/n1464 ) );
  AOI221 U517 ( .A(n575), .B(\position1/N2212 ), .C(n573), .D(n978), .Q(
        \position1/n1268 ) );
  AOI221 U518 ( .A(n542), .B(\position1/N1797 ), .C(n539), .D(n1195), .Q(
        \position1/n1462 ) );
  AOI221 U519 ( .A(n576), .B(\position1/N2214 ), .C(n573), .D(n976), .Q(
        \position1/n1266 ) );
  AOI221 U520 ( .A(n541), .B(\position1/N1791 ), .C(n539), .D(n1201), .Q(
        \position1/n1468 ) );
  AOI221 U521 ( .A(n575), .B(\position1/N2208 ), .C(n573), .D(n982), .Q(
        \position1/n1272 ) );
  AOI221 U522 ( .A(n537), .B(\position1/N1738 ), .C(n535), .D(n1229), .Q(
        \position1/n1494 ) );
  AOI221 U523 ( .A(n571), .B(\position1/N2155 ), .C(n569), .D(n1010), .Q(
        \position1/n1298 ) );
  AOI221 U524 ( .A(n537), .B(\position1/N1740 ), .C(n535), .D(n1226), .Q(
        \position1/n1492 ) );
  AOI221 U525 ( .A(n571), .B(\position1/N2157 ), .C(n569), .D(n1007), .Q(
        \position1/n1296 ) );
  AOI221 U526 ( .A(n537), .B(\position1/N1742 ), .C(n535), .D(n1224), .Q(
        \position1/n1490 ) );
  AOI221 U527 ( .A(n571), .B(\position1/N2159 ), .C(n569), .D(n1005), .Q(
        \position1/n1294 ) );
  AOI221 U528 ( .A(n538), .B(\position1/N1744 ), .C(n535), .D(n1222), .Q(
        \position1/n1488 ) );
  AOI221 U529 ( .A(n572), .B(\position1/N2161 ), .C(n569), .D(n1003), .Q(
        \position1/n1292 ) );
  AOI221 U530 ( .A(n538), .B(\position1/N1746 ), .C(n535), .D(n1220), .Q(
        \position1/n1486 ) );
  AOI221 U531 ( .A(n572), .B(\position1/N2163 ), .C(n569), .D(n1001), .Q(
        \position1/n1290 ) );
  AOI221 U532 ( .A(n537), .B(\position1/N1734 ), .C(n535), .D(n1237), .Q(
        \position1/n1498 ) );
  AOI221 U533 ( .A(n571), .B(\position1/N2151 ), .C(n569), .D(n1018), .Q(
        \position1/n1302 ) );
  AOI221 U534 ( .A(n537), .B(\position1/N1736 ), .C(n535), .D(n1233), .Q(
        \position1/n1496 ) );
  AOI221 U535 ( .A(n571), .B(\position1/N2153 ), .C(n569), .D(n1014), .Q(
        \position1/n1300 ) );
  AOI221 U536 ( .A(n544), .B(\position1/N1836 ), .C(n543), .D(n1180), .Q(
        \position1/n1450 ) );
  AOI221 U537 ( .A(n578), .B(\position1/N2253 ), .C(n577), .D(n961), .Q(
        \position1/n1254 ) );
  AOI221 U538 ( .A(n545), .B(\position1/N1838 ), .C(n543), .D(n1178), .Q(
        \position1/n1448 ) );
  AOI221 U539 ( .A(n579), .B(\position1/N2255 ), .C(n577), .D(n959), .Q(
        \position1/n1252 ) );
  AOI221 U540 ( .A(n545), .B(\position1/N1840 ), .C(n543), .D(n1176), .Q(
        \position1/n1446 ) );
  AOI221 U541 ( .A(n579), .B(\position1/N2257 ), .C(n577), .D(n957), .Q(
        \position1/n1250 ) );
  AOI221 U542 ( .A(n545), .B(\position1/N1846 ), .C(n543), .D(n1170), .Q(
        \position1/n1440 ) );
  AOI221 U543 ( .A(n579), .B(\position1/N2263 ), .C(n577), .D(n951), .Q(
        \position1/n1244 ) );
  AOI221 U544 ( .A(n546), .B(\position1/N1848 ), .C(n543), .D(n1168), .Q(
        \position1/n1438 ) );
  AOI221 U545 ( .A(n580), .B(\position1/N2265 ), .C(n577), .D(n949), .Q(
        \position1/n1242 ) );
  AOI221 U546 ( .A(n1153), .B(n547), .C(\position1/N1888 ), .D(n548), .Q(
        \position1/n1425 ) );
  AOI221 U547 ( .A(n934), .B(n581), .C(\position1/N2305 ), .D(n582), .Q(
        \position1/n1229 ) );
  AOI221 U548 ( .A(n1146), .B(n547), .C(\position1/N1893 ), .D(n549), .Q(
        \position1/n1420 ) );
  AOI221 U549 ( .A(n927), .B(n581), .C(\position1/N2310 ), .D(n583), .Q(
        \position1/n1224 ) );
  NOR31 U550 ( .A(\position1/N1652 ), .B(\position1/N1654 ), .C(
        \position1/N1653 ), .Q(n1970) );
  NOR31 U551 ( .A(\position1/N2069 ), .B(\position1/N2071 ), .C(
        \position1/N2070 ), .Q(n1636) );
  INV3 U552 ( .A(n523), .Q(n522) );
  INV3 U553 ( .A(n557), .Q(n556) );
  INV3 U554 ( .A(\position1/n1521 ), .Q(n1233) );
  AOI221 U555 ( .A(n533), .B(\position1/N1684 ), .C(n531), .D(
        \position1/N1657 ), .Q(\position1/n1521 ) );
  INV3 U556 ( .A(\position1/n1325 ), .Q(n1014) );
  AOI221 U557 ( .A(n567), .B(\position1/N2101 ), .C(n565), .D(
        \position1/N2074 ), .Q(\position1/n1325 ) );
  INV3 U558 ( .A(\position1/n1505 ), .Q(n1214) );
  AOI221 U559 ( .A(n534), .B(\position1/N1700 ), .C(n531), .D(
        \position1/N1673 ), .Q(\position1/n1505 ) );
  XNR21 U560 ( .A(\position1/N1673 ), .B(\position1/sub_216_I4/carry [23]), 
        .Q(\position1/N1700 ) );
  INV3 U561 ( .A(\position1/n1309 ), .Q(n995) );
  AOI221 U562 ( .A(n568), .B(\position1/N2117 ), .C(n565), .D(
        \position1/N2090 ), .Q(\position1/n1309 ) );
  XNR21 U563 ( .A(\position1/N2090 ), .B(\position1/sub_226_I4/carry [23]), 
        .Q(\position1/N2117 ) );
  NOR21 U564 ( .A(\position1/sub_216_I4/carry [23]), .B(\position1/N1673 ), 
        .Q(n115) );
  NOR21 U565 ( .A(\position1/sub_226_I4/carry [23]), .B(\position1/N2090 ), 
        .Q(n131) );
  INV3 U566 ( .A(\position1/n1449 ), .Q(n1152) );
  AOI221 U567 ( .A(n545), .B(\position1/N1837 ), .C(n543), .D(n1179), .Q(
        \position1/n1449 ) );
  INV3 U568 ( .A(\position1/n1253 ), .Q(n933) );
  AOI221 U569 ( .A(n579), .B(\position1/N2254 ), .C(n577), .D(n960), .Q(
        \position1/n1253 ) );
  INV3 U570 ( .A(\position1/n1518 ), .Q(n1228) );
  AOI221 U571 ( .A(n533), .B(\position1/N1687 ), .C(n531), .D(
        \position1/N1660 ), .Q(\position1/n1518 ) );
  INV3 U572 ( .A(\position1/n1322 ), .Q(n1009) );
  AOI221 U573 ( .A(n567), .B(\position1/N2104 ), .C(n565), .D(
        \position1/N2077 ), .Q(\position1/n1322 ) );
  INV3 U574 ( .A(\position1/n1506 ), .Q(n1215) );
  AOI221 U575 ( .A(n534), .B(\position1/N1699 ), .C(n531), .D(
        \position1/N1672 ), .Q(\position1/n1506 ) );
  INV3 U576 ( .A(\position1/n1310 ), .Q(n996) );
  AOI221 U577 ( .A(n568), .B(\position1/N2116 ), .C(n565), .D(
        \position1/N2089 ), .Q(\position1/n1310 ) );
  INV3 U578 ( .A(\position1/n1484 ), .Q(n1191) );
  AOI221 U579 ( .A(n538), .B(\position1/N1748 ), .C(n535), .D(n1218), .Q(
        \position1/n1484 ) );
  INV3 U580 ( .A(\position1/n1288 ), .Q(n972) );
  AOI221 U581 ( .A(n572), .B(\position1/N2165 ), .C(n569), .D(n999), .Q(
        \position1/n1288 ) );
  INV3 U582 ( .A(\position1/N1655 ), .Q(n1264) );
  INV3 U583 ( .A(\position1/N2072 ), .Q(n1045) );
  INV3 U584 ( .A(\position1/n1444 ), .Q(n1144) );
  AOI221 U585 ( .A(n545), .B(\position1/N1842 ), .C(n543), .D(n1174), .Q(
        \position1/n1444 ) );
  INV3 U586 ( .A(\position1/n1248 ), .Q(n925) );
  AOI221 U587 ( .A(n579), .B(\position1/N2259 ), .C(n577), .D(n955), .Q(
        \position1/n1248 ) );
  INV3 U588 ( .A(\position1/n1457 ), .Q(n1162) );
  AOI221 U589 ( .A(n542), .B(\position1/N1802 ), .C(n539), .D(n1188), .Q(
        \position1/n1457 ) );
  XNR21 U590 ( .A(n1188), .B(\position1/sub_216_I6/carry [21]), .Q(
        \position1/N1802 ) );
  INV3 U591 ( .A(\position1/n1261 ), .Q(n943) );
  AOI221 U592 ( .A(n576), .B(\position1/N2219 ), .C(n573), .D(n969), .Q(
        \position1/n1261 ) );
  XNR21 U593 ( .A(n969), .B(\position1/sub_226_I6/carry [21]), .Q(
        \position1/N2219 ) );
  NOR21 U594 ( .A(\position1/N1651 ), .B(\position1/N1677 ), .Q(n1971) );
  NOR21 U595 ( .A(\position1/N2068 ), .B(\position1/N2094 ), .Q(n1637) );
  INV3 U596 ( .A(\position1/n1542 ), .Q(n1288) );
  INV3 U597 ( .A(\position1/n1346 ), .Q(n1069) );
  INV3 U598 ( .A(\position1/n1540 ), .Q(n1284) );
  INV3 U599 ( .A(\position1/n1344 ), .Q(n1065) );
  INV3 U600 ( .A(\position1/n1538 ), .Q(n1280) );
  INV3 U601 ( .A(\position1/n1342 ), .Q(n1061) );
  INV3 U602 ( .A(\position1/n1536 ), .Q(n1276) );
  INV3 U603 ( .A(\position1/n1340 ), .Q(n1057) );
  INV3 U604 ( .A(\position1/n1534 ), .Q(n1272) );
  INV3 U605 ( .A(\position1/n1338 ), .Q(n1053) );
  INV3 U606 ( .A(\position1/n1532 ), .Q(n1268) );
  INV3 U607 ( .A(\position1/n1336 ), .Q(n1049) );
  INV3 U608 ( .A(\position1/n1434 ), .Q(n1130) );
  AOI221 U609 ( .A(n546), .B(\position1/N1852 ), .C(n543), .D(n1164), .Q(
        \position1/n1434 ) );
  INV3 U610 ( .A(\position1/n1238 ), .Q(n911) );
  AOI221 U611 ( .A(n580), .B(\position1/N2269 ), .C(n577), .D(n945), .Q(
        \position1/n1238 ) );
  INV3 U612 ( .A(\position1/n1475 ), .Q(n1180) );
  INV3 U613 ( .A(\position1/n1279 ), .Q(n961) );
  INV3 U614 ( .A(\position1/n1433 ), .Q(n1129) );
  AOI221 U615 ( .A(n546), .B(\position1/N1853 ), .C(n543), .D(n1163), .Q(
        \position1/n1433 ) );
  XNR21 U616 ( .A(n1163), .B(\position1/sub_216_I7/carry [20]), .Q(
        \position1/N1853 ) );
  INV3 U617 ( .A(\position1/n1237 ), .Q(n910) );
  AOI221 U618 ( .A(n580), .B(\position1/N2270 ), .C(n577), .D(n944), .Q(
        \position1/n1237 ) );
  XNR21 U619 ( .A(n944), .B(\position1/sub_226_I7/carry [20]), .Q(
        \position1/N2270 ) );
  INV3 U620 ( .A(\position1/n1481 ), .Q(n1187) );
  AOI221 U621 ( .A(n538), .B(\position1/N1751 ), .C(n535), .D(n1215), .Q(
        \position1/n1481 ) );
  XNR21 U622 ( .A(n1215), .B(\position1/sub_216_I5/carry [22]), .Q(
        \position1/N1751 ) );
  INV3 U623 ( .A(\position1/n1285 ), .Q(n968) );
  AOI221 U624 ( .A(n572), .B(\position1/N2168 ), .C(n569), .D(n996), .Q(
        \position1/n1285 ) );
  XNR21 U625 ( .A(n996), .B(\position1/sub_226_I5/carry [22]), .Q(
        \position1/N2168 ) );
  INV3 U626 ( .A(\position1/n1499 ), .Q(n1207) );
  INV3 U627 ( .A(\position1/n1303 ), .Q(n988) );
  INV3 U628 ( .A(\position1/n1482 ), .Q(n1188) );
  AOI221 U629 ( .A(n538), .B(\position1/N1750 ), .C(n535), .D(n1216), .Q(
        \position1/n1482 ) );
  INV3 U630 ( .A(\position1/n1286 ), .Q(n969) );
  AOI221 U631 ( .A(n572), .B(\position1/N2167 ), .C(n569), .D(n997), .Q(
        \position1/n1286 ) );
  INV3 U632 ( .A(\position1/n1458 ), .Q(n1163) );
  AOI221 U633 ( .A(n542), .B(\position1/N1801 ), .C(n539), .D(n1189), .Q(
        \position1/n1458 ) );
  INV3 U634 ( .A(\position1/n1262 ), .Q(n944) );
  AOI221 U635 ( .A(n576), .B(\position1/N2218 ), .C(n573), .D(n970), .Q(
        \position1/n1262 ) );
  INV3 U636 ( .A(\position1/n1527 ), .Q(n1242) );
  AOI221 U637 ( .A(n532), .B(\position1/N1651 ), .C(n531), .D(
        \position1/N1651 ), .Q(\position1/n1527 ) );
  INV3 U638 ( .A(\position1/n1331 ), .Q(n1023) );
  AOI221 U639 ( .A(n566), .B(\position1/N2068 ), .C(n565), .D(
        \position1/N2068 ), .Q(\position1/n1331 ) );
  INV3 U640 ( .A(\position1/n1528 ), .Q(n1243) );
  AOI221 U641 ( .A(n532), .B(\position1/N1677 ), .C(n531), .D(
        \position1/N1677 ), .Q(\position1/n1528 ) );
  INV3 U642 ( .A(\position1/n1332 ), .Q(n1024) );
  AOI221 U643 ( .A(n566), .B(\position1/N2094 ), .C(n565), .D(
        \position1/N2094 ), .Q(\position1/n1332 ) );
  INV3 U644 ( .A(\position1/n1442 ), .Q(n1142) );
  AOI221 U645 ( .A(n545), .B(\position1/N1844 ), .C(n543), .D(n1172), .Q(
        \position1/n1442 ) );
  INV3 U646 ( .A(\position1/n1246 ), .Q(n923) );
  AOI221 U647 ( .A(n579), .B(\position1/N2261 ), .C(n577), .D(n953), .Q(
        \position1/n1246 ) );
  INV3 U648 ( .A(\position1/n1526 ), .Q(n1241) );
  AOI221 U649 ( .A(n532), .B(\position1/N1652 ), .C(n531), .D(
        \position1/N1652 ), .Q(\position1/n1526 ) );
  INV3 U650 ( .A(\position1/n1330 ), .Q(n1022) );
  AOI221 U651 ( .A(n566), .B(\position1/N2069 ), .C(n565), .D(
        \position1/N2069 ), .Q(\position1/n1330 ) );
  INV3 U652 ( .A(\position1/n1525 ), .Q(n1240) );
  AOI221 U653 ( .A(n532), .B(\position1/N1653 ), .C(n531), .D(
        \position1/N1653 ), .Q(\position1/n1525 ) );
  INV3 U654 ( .A(\position1/n1329 ), .Q(n1021) );
  AOI221 U655 ( .A(n566), .B(\position1/N2070 ), .C(n565), .D(
        \position1/N2070 ), .Q(\position1/n1329 ) );
  INV3 U656 ( .A(\position1/n1504 ), .Q(n1213) );
  AOI221 U657 ( .A(n534), .B(\position1/N1701 ), .C(n531), .D(
        \position1/N1674 ), .Q(\position1/n1504 ) );
  XNR21 U658 ( .A(\position1/sub_216_I4/carry [24]), .B(\position1/N1674 ), 
        .Q(\position1/N1701 ) );
  INV3 U659 ( .A(n115), .Q(\position1/sub_216_I4/carry [24]) );
  INV3 U660 ( .A(\position1/n1308 ), .Q(n994) );
  AOI221 U661 ( .A(n568), .B(\position1/N2118 ), .C(n565), .D(
        \position1/N2091 ), .Q(\position1/n1308 ) );
  XNR21 U662 ( .A(\position1/sub_226_I4/carry [24]), .B(\position1/N2091 ), 
        .Q(\position1/N2118 ) );
  INV3 U663 ( .A(n131), .Q(\position1/sub_226_I4/carry [24]) );
  BUF2 U664 ( .A(\position1/N1883 ), .Q(n548) );
  BUF2 U665 ( .A(\position1/N2300 ), .Q(n582) );
  INV3 U666 ( .A(\position1/n1483 ), .Q(n1189) );
  AOI221 U667 ( .A(n538), .B(\position1/N1749 ), .C(n535), .D(n1217), .Q(
        \position1/n1483 ) );
  INV3 U668 ( .A(\position1/n1287 ), .Q(n970) );
  AOI221 U669 ( .A(n572), .B(\position1/N2166 ), .C(n569), .D(n998), .Q(
        \position1/n1287 ) );
  BUF2 U670 ( .A(\position1/N1831 ), .Q(n544) );
  BUF2 U671 ( .A(\position1/N2248 ), .Q(n578) );
  BUF2 U672 ( .A(\position1/N1675 ), .Q(n532) );
  BUF2 U673 ( .A(\position1/N2092 ), .Q(n566) );
  BUF2 U674 ( .A(\position1/N1727 ), .Q(n536) );
  BUF2 U675 ( .A(\position1/N2144 ), .Q(n570) );
  BUF2 U676 ( .A(\position1/N1779 ), .Q(n540) );
  BUF2 U677 ( .A(\position1/N2196 ), .Q(n574) );
  BUF2 U678 ( .A(\position1/N1831 ), .Q(n545) );
  BUF2 U679 ( .A(\position1/N2248 ), .Q(n579) );
  BUF2 U680 ( .A(\position1/N1675 ), .Q(n533) );
  BUF2 U681 ( .A(\position1/N2092 ), .Q(n567) );
  BUF2 U682 ( .A(\position1/N1727 ), .Q(n537) );
  BUF2 U683 ( .A(\position1/N2144 ), .Q(n571) );
  BUF2 U684 ( .A(\position1/N1779 ), .Q(n541) );
  BUF2 U685 ( .A(\position1/N2196 ), .Q(n575) );
  BUF2 U686 ( .A(n530), .Q(n528) );
  INV3 U687 ( .A(\position1/N1623 ), .Q(n530) );
  BUF2 U688 ( .A(n564), .Q(n562) );
  INV3 U689 ( .A(\position1/N2040 ), .Q(n564) );
  BUF2 U690 ( .A(\position1/N1883 ), .Q(n549) );
  BUF2 U691 ( .A(\position1/N2300 ), .Q(n583) );
  BUF2 U692 ( .A(\position1/N1883 ), .Q(n550) );
  BUF2 U693 ( .A(\position1/N2300 ), .Q(n584) );
  BUF2 U694 ( .A(\position1/N1831 ), .Q(n546) );
  BUF2 U695 ( .A(\position1/N2248 ), .Q(n580) );
  BUF2 U696 ( .A(\position1/N1675 ), .Q(n534) );
  BUF2 U697 ( .A(\position1/N2092 ), .Q(n568) );
  BUF2 U698 ( .A(\position1/N1727 ), .Q(n538) );
  BUF2 U699 ( .A(\position1/N2144 ), .Q(n572) );
  BUF2 U700 ( .A(\position1/N1779 ), .Q(n542) );
  BUF2 U701 ( .A(\position1/N2196 ), .Q(n576) );
  INV3 U702 ( .A(n116), .Q(\position1/sub_216_I5/carry [23]) );
  NOR21 U703 ( .A(\position1/sub_216_I5/carry [22]), .B(n1215), .Q(n116) );
  INV3 U704 ( .A(n132), .Q(\position1/sub_226_I5/carry [23]) );
  NOR21 U705 ( .A(\position1/sub_226_I5/carry [22]), .B(n996), .Q(n132) );
  INV3 U706 ( .A(n118), .Q(\position1/sub_216_I6/carry [22]) );
  NOR21 U707 ( .A(\position1/sub_216_I6/carry [21]), .B(n1188), .Q(n118) );
  INV3 U708 ( .A(n134), .Q(\position1/sub_226_I6/carry [22]) );
  NOR21 U709 ( .A(\position1/sub_226_I6/carry [21]), .B(n969), .Q(n134) );
  INV3 U710 ( .A(n121), .Q(\position1/sub_216_I7/carry [21]) );
  NOR21 U711 ( .A(\position1/sub_216_I7/carry [20]), .B(n1163), .Q(n121) );
  INV3 U712 ( .A(n125), .Q(\position1/sub_216_I8/carry [20]) );
  NOR21 U713 ( .A(\position1/sub_216_I8/carry [19]), .B(n1130), .Q(n125) );
  INV3 U714 ( .A(n137), .Q(\position1/sub_226_I7/carry [21]) );
  NOR21 U715 ( .A(\position1/sub_226_I7/carry [20]), .B(n944), .Q(n137) );
  INV3 U716 ( .A(n141), .Q(\position1/sub_226_I8/carry [20]) );
  NOR21 U717 ( .A(\position1/sub_226_I8/carry [19]), .B(n911), .Q(n141) );
  NOR21 U718 ( .A(n1144), .B(n40), .Q(n1841) );
  NOR21 U719 ( .A(n925), .B(n40), .Q(n1507) );
  NAND22 U720 ( .A(n1167), .B(n42), .Q(n1885) );
  NAND22 U721 ( .A(n948), .B(n42), .Q(n1551) );
  INV3 U722 ( .A(\position1/n1418 ), .Q(n1112) );
  AOI221 U723 ( .A(n1143), .B(n547), .C(\position1/N1895 ), .D(n549), .Q(
        \position1/n1418 ) );
  INV3 U724 ( .A(\position1/n1222 ), .Q(n893) );
  AOI221 U725 ( .A(n924), .B(n581), .C(\position1/N2312 ), .D(n583), .Q(
        \position1/n1222 ) );
  INV3 U726 ( .A(\position1/n1409 ), .Q(n1103) );
  AOI221 U727 ( .A(n1130), .B(n547), .C(\position1/N1904 ), .D(n550), .Q(
        \position1/n1409 ) );
  XNR21 U728 ( .A(n1130), .B(\position1/sub_216_I8/carry [19]), .Q(
        \position1/N1904 ) );
  INV3 U729 ( .A(\position1/n1213 ), .Q(n884) );
  AOI221 U730 ( .A(n911), .B(n581), .C(\position1/N2321 ), .D(n584), .Q(
        \position1/n1213 ) );
  XNR21 U731 ( .A(n911), .B(\position1/sub_226_I8/carry [19]), .Q(
        \position1/N2321 ) );
  INV3 U732 ( .A(\position1/n1410 ), .Q(n1104) );
  AOI221 U733 ( .A(n1132), .B(n547), .C(\position1/N1903 ), .D(n550), .Q(
        \position1/n1410 ) );
  INV3 U734 ( .A(\position1/n1214 ), .Q(n885) );
  AOI221 U735 ( .A(n913), .B(n581), .C(\position1/N2320 ), .D(n584), .Q(
        \position1/n1214 ) );
  BUF2 U736 ( .A(\position1/N1883 ), .Q(n551) );
  BUF2 U737 ( .A(\position1/N2300 ), .Q(n585) );
  INV3 U738 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[0] ), .Q(
        n809) );
  NAND22 U739 ( .A(cam_y[0]), .B(n1361), .Q(
        \position1/dp_cluster_5/mult_add_179_aco/PROD_not[0] ) );
  INV3 U740 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[0] ), .Q(
        n852) );
  NAND22 U741 ( .A(cam_x[0]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[0] ) );
  INV3 U742 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[0] ), .Q(
        n853) );
  NAND22 U743 ( .A(cam_x[0]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[0] ) );
  BUF2 U744 ( .A(n2130), .Q(cam_x[4]) );
  INV3 U745 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[0] ), .Q(
        n810) );
  NAND22 U746 ( .A(cam_y[0]), .B(n1360), .Q(
        \position1/dp_cluster_1/mult_add_197_aco/PROD_not[0] ) );
  BUF2 U747 ( .A(n2130), .Q(n495) );
  BUF2 U748 ( .A(n2128), .Q(cam_x[6]) );
  BUF2 U749 ( .A(n2128), .Q(n491) );
  AOI221 U750 ( .A(\position1/N606 ), .B(n479), .C(\position1/N577 ), .D(n478), 
        .Q(\position1/n1068 ) );
  XOR21 U751 ( .A(n586), .B(\position1/r458/carry [17]), .Q(\position1/N577 )
         );
  XOR21 U752 ( .A(\position1/r416/carry [17]), .B(n586), .Q(\position1/N606 )
         );
  NOR21 U753 ( .A(n300), .B(n301), .Q(\position1/r458/carry [17]) );
  INV3 U754 ( .A(\position1/n1066 ), .Q(n672) );
  AOI221 U755 ( .A(n633), .B(n586), .C(\position1/n1067 ), .D(n741), .Q(
        \position1/n1066 ) );
  NAND22 U756 ( .A(\position1/n1068 ), .B(\position1/n1069 ), .Q(
        \position1/n1067 ) );
  AOI221 U757 ( .A(n2), .B(n477), .C(\position1/N447 ), .D(n476), .Q(
        \position1/n1069 ) );
  XNR21 U758 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .B(
        \position1/sub_250_3/carry[5] ), .Q(\position1/N2387 ) );
  XNR21 U759 ( .A(n493), .B(\position1/sub_250/carry[5] ), .Q(
        \position1/N2377 ) );
  XNR21 U760 ( .A(n489), .B(\position1/sub_250/carry[7] ), .Q(
        \position1/N2379 ) );
  NOR21 U761 ( .A(\position1/n1056 ), .B(\position1/n1057 ), .Q(
        \position1/n856 ) );
  XOR21 U762 ( .A(cam_x[2]), .B(\position1/sub_250/carry[2] ), .Q(
        \position1/N2374 ) );
  XOR21 U763 ( .A(n497), .B(\position1/add_250/carry[3] ), .Q(
        \position1/N2396 ) );
  XOR21 U764 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .B(
        \position1/add_250_2/carry[5] ), .Q(\position1/N2409 ) );
  XOR21 U765 ( .A(n493), .B(\position1/add_250/carry[5] ), .Q(
        \position1/N2398 ) );
  XOR21 U766 ( .A(n489), .B(\position1/add_250/carry[7] ), .Q(
        \position1/N2400 ) );
  XNR21 U767 ( .A(cam_x[3]), .B(\position1/sub_250/carry[3] ), .Q(
        \position1/N2375 ) );
  XNR21 U768 ( .A(n499), .B(\position1/add_250/carry[2] ), .Q(
        \position1/N2395 ) );
  BUF2 U769 ( .A(\position1/n857 ), .Q(n640) );
  BUF2 U770 ( .A(\position1/n857 ), .Q(n639) );
  AOI221 U771 ( .A(\position1/N537 ), .B(n512), .C(\position1/N981 ), .D(n640), 
        .Q(\position1/n946 ) );
  AOI221 U772 ( .A(\position1/N538 ), .B(n512), .C(\position1/N982 ), .D(n640), 
        .Q(\position1/n942 ) );
  AOI221 U773 ( .A(\position1/N539 ), .B(n740), .C(\position1/N983 ), .D(n640), 
        .Q(\position1/n938 ) );
  AOI221 U774 ( .A(\position1/N540 ), .B(n511), .C(\position1/N984 ), .D(n640), 
        .Q(\position1/n934 ) );
  AOI221 U775 ( .A(\position1/N487 ), .B(n740), .C(\position1/N906 ), .D(n641), 
        .Q(\position1/n1046 ) );
  AOI221 U776 ( .A(\position1/N488 ), .B(n740), .C(\position1/N907 ), .D(n641), 
        .Q(\position1/n1042 ) );
  AOI221 U777 ( .A(\position1/N489 ), .B(n740), .C(\position1/N908 ), .D(n640), 
        .Q(\position1/n1038 ) );
  NOR21 U778 ( .A(n303), .B(n304), .Q(\position1/sub_250/carry[3] ) );
  INV3 U779 ( .A(cam_x[2]), .Q(n304) );
  INV3 U780 ( .A(\position1/sub_250/carry[2] ), .Q(n303) );
  INV3 U781 ( .A(\position1/n1179 ), .Q(n712) );
  BUF2 U782 ( .A(\position1/n857 ), .Q(n641) );
  INV3 U783 ( .A(\position1/n1059 ), .Q(n740) );
  NAND22 U784 ( .A(n741), .B(n478), .Q(\position1/n1059 ) );
  INV3 U785 ( .A(\position1/n1141 ), .Q(n782) );
  INV3 U786 ( .A(n147), .Q(\position1/sub_250/carry[4] ) );
  NOR21 U787 ( .A(\position1/sub_250/carry[3] ), .B(cam_x[3]), .Q(n147) );
  INV3 U788 ( .A(n157), .Q(\position1/add_250/carry[2] ) );
  NOR21 U789 ( .A(cam_x[0]), .B(n501), .Q(n157) );
  INV3 U790 ( .A(n149), .Q(\position1/sub_250/carry[6] ) );
  NOR21 U791 ( .A(\position1/sub_250/carry[5] ), .B(n493), .Q(n149) );
  INV3 U792 ( .A(n154), .Q(\position1/sub_250_3/carry[6] ) );
  NOR21 U793 ( .A(\position1/sub_250_3/carry[5] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), .Q(n154) );
  INV3 U794 ( .A(n158), .Q(\position1/add_250/carry[3] ) );
  NOR21 U795 ( .A(\position1/add_250/carry[2] ), .B(n499), .Q(n158) );
  INV3 U796 ( .A(\position1/N2408 ), .Q(n797) );
  INV3 U797 ( .A(\position1/N2410 ), .Q(n789) );
  INV3 U798 ( .A(\position1/N2412 ), .Q(n779) );
  INV3 U799 ( .A(\position1/N2401 ), .Q(n836) );
  INV3 U800 ( .A(\position1/N2411 ), .Q(n785) );
  INV3 U801 ( .A(\position1/N2380 ), .Q(n844) );
  NOR21 U802 ( .A(cam_x[1]), .B(n503), .Q(\position1/n1399 ) );
  NOR40 U803 ( .A(n864), .B(\position1/n1398 ), .C(cam_x[5]), .D(cam_x[4]), 
        .Q(\position1/n1397 ) );
  AOI221 U804 ( .A(\position1/n1399 ), .B(cam_x[2]), .C(cam_x[0]), .D(n304), 
        .Q(\position1/n1398 ) );
  INV3 U805 ( .A(\position1/n1400 ), .Q(n864) );
  NOR21 U806 ( .A(n211), .B(n302), .Q(\position1/sub_250/carry[2] ) );
  INV3 U807 ( .A(n501), .Q(n302) );
  NOR21 U808 ( .A(n309), .B(n310), .Q(\position1/add_250/carry[6] ) );
  INV3 U809 ( .A(n493), .Q(n310) );
  INV3 U810 ( .A(\position1/add_250/carry[5] ), .Q(n309) );
  NOR21 U811 ( .A(n316), .B(\gensync1/n94 ), .Q(\position1/add_250_2/carry[6] ) );
  INV3 U812 ( .A(\position1/add_250_2/carry[5] ), .Q(n316) );
  NOR21 U813 ( .A(n158), .B(n306), .Q(\position1/add_250/carry[4] ) );
  INV3 U814 ( .A(n497), .Q(n306) );
  NOR21 U815 ( .A(\position1/n1063 ), .B(\position1/n1064 ), .Q(
        \position1/n859 ) );
  BUF2 U816 ( .A(n673), .Q(n509) );
  BUF2 U817 ( .A(n673), .Q(n508) );
  BUF2 U818 ( .A(\position1/n858 ), .Q(n643) );
  BUF2 U819 ( .A(\position1/n858 ), .Q(n642) );
  BUF2 U820 ( .A(\position1/n858 ), .Q(n644) );
  BUF2 U821 ( .A(n673), .Q(n510) );
  INV3 U822 ( .A(\gensync1/n103 ), .Q(IMG_top) );
  INV3 U823 ( .A(\position1/r458/carry [16]), .Q(n301) );
  NOR21 U824 ( .A(\position1/n1064 ), .B(n482), .Q(n480) );
  NOR21 U825 ( .A(\position1/n1064 ), .B(n482), .Q(n481) );
  NOR21 U826 ( .A(\position1/n1064 ), .B(n482), .Q(\position1/n1154 ) );
  NAND22 U827 ( .A(\image_process1/n57 ), .B(n876), .Q(\image_process1/n97 )
         );
  INV3 U828 ( .A(\position1/n1064 ), .Q(n741) );
  BUF2 U829 ( .A(\position1/n834 ), .Q(n633) );
  INV3 U830 ( .A(\position1/n1056 ), .Q(n1359) );
  INV3 U831 ( .A(n587), .Q(n586) );
  NAND22 U832 ( .A(\image_process1/n113 ), .B(n876), .Q(\image_process1/n56 )
         );
  BUF2 U833 ( .A(\position1/n834 ), .Q(n634) );
  INV3 U834 ( .A(n2043), .Q(n1265) );
  AOI211 U835 ( .A(n2044), .B(n2), .C(\position1/n1530 ), .Q(n2043) );
  AOI221 U836 ( .A(n2042), .B(n2041), .C(n44), .D(n1267), .Q(n2044) );
  INV3 U837 ( .A(n1709), .Q(n1046) );
  AOI211 U838 ( .A(n1710), .B(n2), .C(\position1/n1334 ), .Q(n1709) );
  AOI221 U839 ( .A(n1708), .B(n1707), .C(n44), .D(n1048), .Q(n1710) );
  INV3 U840 ( .A(\position1/N1632 ), .Q(n1297) );
  INV3 U841 ( .A(\position1/N2049 ), .Q(n1078) );
  XOR21 U842 ( .A(n1299), .B(n34), .Q(n104) );
  XOR21 U843 ( .A(n1080), .B(n34), .Q(n105) );
  INV3 U844 ( .A(\position1/N1633 ), .Q(n1294) );
  INV3 U845 ( .A(\position1/N2050 ), .Q(n1075) );
  INV3 U846 ( .A(\position1/N1637 ), .Q(n1285) );
  INV3 U847 ( .A(\position1/N2054 ), .Q(n1066) );
  INV3 U848 ( .A(\position1/N1639 ), .Q(n1281) );
  INV3 U849 ( .A(\position1/N2056 ), .Q(n1062) );
  INV3 U850 ( .A(\position1/N1641 ), .Q(n1277) );
  INV3 U851 ( .A(\position1/N2058 ), .Q(n1058) );
  INV3 U852 ( .A(\position1/N1643 ), .Q(n1273) );
  INV3 U853 ( .A(\position1/N2060 ), .Q(n1054) );
  INV3 U854 ( .A(\position1/N1645 ), .Q(n1269) );
  INV3 U855 ( .A(\position1/N2062 ), .Q(n1050) );
  INV3 U856 ( .A(\position1/N1635 ), .Q(n1289) );
  INV3 U857 ( .A(\position1/N2052 ), .Q(n1070) );
  AOI221 U858 ( .A(n524), .B(\position1/N1582 ), .C(n522), .D(
        \position1/N1555 ), .Q(\position1/n1544 ) );
  AOI221 U859 ( .A(n558), .B(\position1/N1999 ), .C(n556), .D(
        \position1/N1972 ), .Q(\position1/n1348 ) );
  XNR21 U860 ( .A(\position1/sub_216_I3/carry [24]), .B(\position1/n1529 ), 
        .Q(n106) );
  XNR21 U861 ( .A(\position1/sub_226_I3/carry [24]), .B(\position1/n1333 ), 
        .Q(n107) );
  OAI2111 U862 ( .A(n2), .B(\position1/n1459 ), .C(n1894), .D(n1893), .Q(
        \position1/N1831 ) );
  AOI311 U863 ( .A(n1892), .B(n1891), .C(n1890), .D(n1163), .Q(n1894) );
  NOR40 U864 ( .A(n1159), .B(n1160), .C(n1161), .D(n1162), .Q(n1893) );
  NAND22 U865 ( .A(n586), .B(\position1/n1459 ), .Q(n1890) );
  OAI2111 U866 ( .A(n2), .B(\position1/n1263 ), .C(n1560), .D(n1559), .Q(
        \position1/N2248 ) );
  AOI311 U867 ( .A(n1558), .B(n1557), .C(n1556), .D(n944), .Q(n1560) );
  NOR40 U868 ( .A(n940), .B(n941), .C(n942), .D(n943), .Q(n1559) );
  NAND22 U869 ( .A(n586), .B(\position1/n1263 ), .Q(n1556) );
  OAI2111 U870 ( .A(n2), .B(n1244), .C(n2007), .D(n2006), .Q(\position1/N1675 ) );
  INV3 U871 ( .A(n2005), .Q(n1244) );
  NOR21 U872 ( .A(\position1/N1674 ), .B(\position1/N1673 ), .Q(n2006) );
  OAI2111 U873 ( .A(n2), .B(n1025), .C(n1673), .D(n1672), .Q(\position1/N2092 ) );
  INV3 U874 ( .A(n1671), .Q(n1025) );
  NOR21 U875 ( .A(\position1/N2091 ), .B(\position1/N2090 ), .Q(n1672) );
  OAI2111 U876 ( .A(n2), .B(n1969), .C(n1212), .D(n1968), .Q(\position1/N1727 ) );
  INV3 U877 ( .A(n1967), .Q(n1212) );
  NOR31 U878 ( .A(n1215), .B(n1213), .C(n1214), .Q(n1968) );
  AOI211 U879 ( .A(n1969), .B(n2), .C(\position1/n1507 ), .Q(n1967) );
  OAI2111 U880 ( .A(n2), .B(n1635), .C(n993), .D(n1634), .Q(\position1/N2144 )
         );
  INV3 U881 ( .A(n1633), .Q(n993) );
  NOR31 U882 ( .A(n996), .B(n994), .C(n995), .Q(n1634) );
  AOI211 U883 ( .A(n1635), .B(n2), .C(\position1/n1311 ), .Q(n1633) );
  OAI2111 U884 ( .A(n2), .B(n1932), .C(n1931), .D(n1930), .Q(\position1/N1779 ) );
  AOI211 U885 ( .A(n1189), .B(n1929), .C(n1188), .Q(n1931) );
  NOR31 U886 ( .A(n1187), .B(n1185), .C(n1186), .Q(n1930) );
  NAND22 U887 ( .A(n586), .B(n1932), .Q(n1929) );
  OAI2111 U888 ( .A(n2), .B(n1598), .C(n1597), .D(n1596), .Q(\position1/N2196 ) );
  AOI211 U889 ( .A(n970), .B(n1595), .C(n969), .Q(n1597) );
  NOR31 U890 ( .A(n968), .B(n966), .C(n967), .Q(n1596) );
  NAND22 U891 ( .A(n586), .B(n1598), .Q(n1595) );
  INV3 U892 ( .A(\position1/N1647 ), .Q(n1246) );
  INV3 U893 ( .A(\position1/N2064 ), .Q(n1027) );
  AOI221 U894 ( .A(n525), .B(\position1/N1596 ), .C(n522), .D(
        \position1/N1569 ), .Q(\position1/n1530 ) );
  AOI221 U895 ( .A(n559), .B(\position1/N2013 ), .C(n556), .D(
        \position1/N1986 ), .Q(\position1/n1334 ) );
  AOI221 U896 ( .A(n524), .B(\position1/N1584 ), .C(n522), .D(
        \position1/N1557 ), .Q(\position1/n1542 ) );
  AOI221 U897 ( .A(n558), .B(\position1/N2001 ), .C(n556), .D(
        \position1/N1974 ), .Q(\position1/n1346 ) );
  AOI221 U898 ( .A(n524), .B(\position1/N1586 ), .C(n522), .D(
        \position1/N1559 ), .Q(\position1/n1540 ) );
  AOI221 U899 ( .A(n558), .B(\position1/N2003 ), .C(n556), .D(
        \position1/N1976 ), .Q(\position1/n1344 ) );
  AOI221 U900 ( .A(n525), .B(\position1/N1588 ), .C(n522), .D(
        \position1/N1561 ), .Q(\position1/n1538 ) );
  AOI221 U901 ( .A(n559), .B(\position1/N2005 ), .C(n556), .D(
        \position1/N1978 ), .Q(\position1/n1342 ) );
  AOI221 U902 ( .A(n525), .B(\position1/N1590 ), .C(n522), .D(
        \position1/N1563 ), .Q(\position1/n1536 ) );
  AOI221 U903 ( .A(n559), .B(\position1/N2007 ), .C(n556), .D(
        \position1/N1980 ), .Q(\position1/n1340 ) );
  AOI221 U904 ( .A(n525), .B(\position1/N1592 ), .C(n522), .D(
        \position1/N1565 ), .Q(\position1/n1534 ) );
  AOI221 U905 ( .A(n559), .B(\position1/N2009 ), .C(n556), .D(
        \position1/N1982 ), .Q(\position1/n1338 ) );
  AOI221 U906 ( .A(n525), .B(\position1/N1594 ), .C(n522), .D(
        \position1/N1567 ), .Q(\position1/n1532 ) );
  AOI221 U907 ( .A(n559), .B(\position1/N2011 ), .C(n556), .D(
        \position1/N1984 ), .Q(\position1/n1336 ) );
  AOI221 U908 ( .A(n537), .B(\position1/N1733 ), .C(n535), .D(n1239), .Q(
        \position1/n1499 ) );
  XNR21 U909 ( .A(n1239), .B(n34), .Q(\position1/N1733 ) );
  AOI221 U910 ( .A(n571), .B(\position1/N2150 ), .C(n569), .D(n1020), .Q(
        \position1/n1303 ) );
  XNR21 U911 ( .A(n1020), .B(n34), .Q(\position1/N2150 ) );
  AOI221 U912 ( .A(n540), .B(\position1/N1784 ), .C(n539), .D(n1208), .Q(
        \position1/n1475 ) );
  XNR21 U913 ( .A(n1208), .B(n34), .Q(\position1/N1784 ) );
  AOI221 U914 ( .A(n574), .B(\position1/N2201 ), .C(n573), .D(n989), .Q(
        \position1/n1279 ) );
  XNR21 U915 ( .A(n989), .B(n34), .Q(\position1/N2201 ) );
  NAND22 U916 ( .A(n1857), .B(n1856), .Q(\position1/N1883 ) );
  NOR40 U917 ( .A(n1129), .B(n1130), .C(n1855), .D(n1854), .Q(n1857) );
  NOR40 U918 ( .A(n1125), .B(n1126), .C(n1127), .D(n1128), .Q(n1856) );
  NOR21 U919 ( .A(n586), .B(\position1/n1435 ), .Q(n1854) );
  NAND22 U920 ( .A(n1523), .B(n1522), .Q(\position1/N2300 ) );
  NOR40 U921 ( .A(n910), .B(n911), .C(n1521), .D(n1520), .Q(n1523) );
  NOR40 U922 ( .A(n906), .B(n907), .C(n908), .D(n909), .Q(n1522) );
  NOR21 U923 ( .A(n586), .B(\position1/n1239 ), .Q(n1520) );
  INV3 U924 ( .A(n521), .Q(n520) );
  INV3 U925 ( .A(n555), .Q(n554) );
  INV3 U926 ( .A(n521), .Q(n519) );
  INV3 U927 ( .A(n555), .Q(n553) );
  INV3 U928 ( .A(n521), .Q(n518) );
  INV3 U929 ( .A(n555), .Q(n552) );
  INV3 U930 ( .A(\position1/n1523 ), .Q(n1237) );
  AOI221 U931 ( .A(n533), .B(\position1/N1682 ), .C(n531), .D(
        \position1/N1655 ), .Q(\position1/n1523 ) );
  XNR21 U932 ( .A(\position1/N1655 ), .B(n34), .Q(\position1/N1682 ) );
  INV3 U933 ( .A(\position1/n1327 ), .Q(n1018) );
  AOI221 U934 ( .A(n567), .B(\position1/N2099 ), .C(n565), .D(
        \position1/N2072 ), .Q(\position1/n1327 ) );
  XNR21 U935 ( .A(\position1/N2072 ), .B(n513), .Q(\position1/N2099 ) );
  INV3 U936 ( .A(\position1/n1451 ), .Q(n1155) );
  AOI221 U937 ( .A(n544), .B(\position1/N1835 ), .C(n543), .D(n1181), .Q(
        \position1/n1451 ) );
  XNR21 U938 ( .A(n1181), .B(n513), .Q(\position1/N1835 ) );
  INV3 U939 ( .A(\position1/n1255 ), .Q(n936) );
  AOI221 U940 ( .A(n578), .B(\position1/N2252 ), .C(n577), .D(n962), .Q(
        \position1/n1255 ) );
  XNR21 U941 ( .A(n962), .B(n34), .Q(\position1/N2252 ) );
  INV3 U942 ( .A(\position1/n1547 ), .Q(n1299) );
  INV3 U943 ( .A(\position1/n1351 ), .Q(n1080) );
  NAND31 U944 ( .A(\position1/n1550 ), .B(\position1/n1548 ), .C(
        \position1/n1549 ), .Q(n108) );
  NAND31 U945 ( .A(\position1/n1354 ), .B(\position1/n1352 ), .C(
        \position1/n1353 ), .Q(n109) );
  INV3 U946 ( .A(\position1/n1543 ), .Q(n1291) );
  INV3 U947 ( .A(\position1/n1347 ), .Q(n1072) );
  INV3 U948 ( .A(\position1/n1546 ), .Q(n1298) );
  INV3 U949 ( .A(\position1/n1350 ), .Q(n1079) );
  INV3 U950 ( .A(\position1/n1541 ), .Q(n1286) );
  INV3 U951 ( .A(\position1/n1345 ), .Q(n1067) );
  INV3 U952 ( .A(\position1/n1539 ), .Q(n1282) );
  INV3 U953 ( .A(\position1/n1343 ), .Q(n1063) );
  INV3 U954 ( .A(\position1/n1537 ), .Q(n1278) );
  INV3 U955 ( .A(\position1/n1341 ), .Q(n1059) );
  INV3 U956 ( .A(\position1/n1535 ), .Q(n1274) );
  INV3 U957 ( .A(\position1/n1339 ), .Q(n1055) );
  INV3 U958 ( .A(\position1/N1569 ), .Q(n1301) );
  INV3 U959 ( .A(\position1/N1986 ), .Q(n1082) );
  INV3 U960 ( .A(\position1/n1533 ), .Q(n1270) );
  INV3 U961 ( .A(\position1/n1337 ), .Q(n1051) );
  INV3 U962 ( .A(\position1/n1531 ), .Q(n1267) );
  INV3 U963 ( .A(\position1/n1335 ), .Q(n1048) );
  INV3 U964 ( .A(\position1/n1334 ), .Q(n1047) );
  INV3 U965 ( .A(\position1/n1530 ), .Q(n1266) );
  INV3 U966 ( .A(n167), .Q(\position1/sub_216_I3/carry [7]) );
  NOR21 U967 ( .A(n513), .B(n1299), .Q(n167) );
  INV3 U968 ( .A(n173), .Q(\position1/sub_226_I3/carry [7]) );
  NOR21 U969 ( .A(n513), .B(n1080), .Q(n173) );
  INV3 U970 ( .A(\position1/n1545 ), .Q(n1296) );
  INV3 U971 ( .A(\position1/n1349 ), .Q(n1077) );
  INV3 U972 ( .A(\position1/n1544 ), .Q(n1293) );
  INV3 U973 ( .A(\position1/n1348 ), .Q(n1074) );
  INV3 U974 ( .A(n168), .Q(\position1/sub_216_I4/carry [6]) );
  NOR21 U975 ( .A(n513), .B(\position1/N1655 ), .Q(n168) );
  INV3 U976 ( .A(n174), .Q(\position1/sub_226_I4/carry [6]) );
  NOR21 U977 ( .A(n513), .B(\position1/N2072 ), .Q(n174) );
  INV3 U978 ( .A(n169), .Q(\position1/sub_216_I5/carry [5]) );
  NOR21 U979 ( .A(n513), .B(n1239), .Q(n169) );
  INV3 U980 ( .A(n175), .Q(\position1/sub_226_I5/carry [5]) );
  NOR21 U981 ( .A(n34), .B(n1020), .Q(n175) );
  INV3 U982 ( .A(n170), .Q(\position1/sub_216_I6/carry [4]) );
  NOR21 U983 ( .A(n513), .B(n1208), .Q(n170) );
  INV3 U984 ( .A(n171), .Q(\position1/sub_216_I7/carry [3]) );
  NOR21 U985 ( .A(n513), .B(n1181), .Q(n171) );
  INV3 U986 ( .A(n177), .Q(\position1/sub_226_I7/carry [3]) );
  NOR21 U987 ( .A(n34), .B(n962), .Q(n177) );
  INV3 U988 ( .A(n176), .Q(\position1/sub_226_I6/carry [4]) );
  NOR21 U989 ( .A(n34), .B(n989), .Q(n176) );
  INV3 U990 ( .A(n130), .Q(\position1/sub_216_I8/carry [2]) );
  NOR21 U991 ( .A(n513), .B(n1157), .Q(n130) );
  INV3 U992 ( .A(n146), .Q(\position1/sub_226_I8/carry [2]) );
  NOR21 U993 ( .A(n34), .B(n938), .Q(n146) );
  NAND31 U994 ( .A(\position1/n1553 ), .B(\position1/n1551 ), .C(
        \position1/n1552 ), .Q(n110) );
  NAND31 U995 ( .A(\position1/n1357 ), .B(\position1/n1355 ), .C(
        \position1/n1356 ), .Q(n111) );
  AOI221 U996 ( .A(n1157), .B(n547), .C(\position1/N1886 ), .D(n548), .Q(
        \position1/n1427 ) );
  XNR21 U997 ( .A(n1157), .B(n513), .Q(\position1/N1886 ) );
  AOI221 U998 ( .A(n938), .B(n581), .C(\position1/N2303 ), .D(n582), .Q(
        \position1/n1231 ) );
  XNR21 U999 ( .A(n938), .B(n34), .Q(\position1/N2303 ) );
  BUF2 U1000 ( .A(\position1/N1571 ), .Q(n523) );
  BUF2 U1001 ( .A(\position1/N1988 ), .Q(n557) );
  BUF2 U1002 ( .A(\position1/N1571 ), .Q(n524) );
  BUF2 U1003 ( .A(\position1/N1988 ), .Q(n558) );
  MAJ31 U1004 ( .A(\position1/n1411 ), .B(n1815), .C(n2), .Q(n1819) );
  AOI221 U1005 ( .A(n1105), .B(n300), .C(n1814), .D(n1813), .Q(n1815) );
  AOI221 U1006 ( .A(n1133), .B(n547), .C(\position1/N1902 ), .D(n550), .Q(
        \position1/n1411 ) );
  INV3 U1007 ( .A(\position1/n1412 ), .Q(n1105) );
  MAJ31 U1008 ( .A(\position1/n1215 ), .B(n1481), .C(n2), .Q(n1485) );
  AOI221 U1009 ( .A(n886), .B(n300), .C(n1480), .D(n1479), .Q(n1481) );
  AOI221 U1010 ( .A(n914), .B(n581), .C(\position1/N2319 ), .D(n584), .Q(
        \position1/n1215 ) );
  INV3 U1011 ( .A(\position1/n1216 ), .Q(n886) );
  BUF2 U1012 ( .A(\position1/N1571 ), .Q(n525) );
  BUF2 U1013 ( .A(\position1/N1988 ), .Q(n559) );
  NOR21 U1014 ( .A(n1155), .B(n628), .Q(n1826) );
  NOR21 U1015 ( .A(n936), .B(n273), .Q(n1492) );
  NOR21 U1016 ( .A(n1152), .B(n246), .Q(n1825) );
  NOR21 U1017 ( .A(n933), .B(n246), .Q(n1491) );
  NOR21 U1018 ( .A(n1149), .B(n278), .Q(n1824) );
  NOR21 U1019 ( .A(n930), .B(n250), .Q(n1490) );
  NOR21 U1020 ( .A(n1140), .B(n261), .Q(n1823) );
  NOR21 U1021 ( .A(n921), .B(n290), .Q(n1489) );
  NOR21 U1022 ( .A(n1137), .B(n294), .Q(n1822) );
  NOR21 U1023 ( .A(n918), .B(n265), .Q(n1488) );
  NOR21 U1024 ( .A(n1134), .B(n269), .Q(n1821) );
  NOR21 U1025 ( .A(n915), .B(n298), .Q(n1487) );
  NOR21 U1026 ( .A(n485), .B(n547), .Q(\position1/N2355 ) );
  NOR21 U1027 ( .A(n486), .B(n581), .Q(\position1/N2364 ) );
  NOR21 U1028 ( .A(n487), .B(n522), .Q(\position1/N2361 ) );
  NOR21 U1029 ( .A(n486), .B(n556), .Q(\position1/N2370 ) );
  NOR21 U1030 ( .A(n485), .B(n531), .Q(\position1/N2359 ) );
  NOR21 U1031 ( .A(n485), .B(n543), .Q(\position1/N2356 ) );
  NOR21 U1032 ( .A(n487), .B(n577), .Q(\position1/N2365 ) );
  NOR21 U1033 ( .A(n485), .B(n535), .Q(\position1/N2358 ) );
  NOR21 U1034 ( .A(n485), .B(n539), .Q(\position1/N2357 ) );
  NOR21 U1035 ( .A(n486), .B(n565), .Q(\position1/N2368 ) );
  NOR21 U1036 ( .A(n487), .B(n569), .Q(\position1/N2367 ) );
  NOR21 U1037 ( .A(n486), .B(n573), .Q(\position1/N2366 ) );
  INV3 U1038 ( .A(n1827), .Q(n1156) );
  AOI211 U1039 ( .A(n1158), .B(n34), .C(n1157), .Q(n1827) );
  INV3 U1040 ( .A(n1493), .Q(n937) );
  AOI211 U1041 ( .A(n939), .B(n34), .C(n938), .Q(n1493) );
  NOR21 U1042 ( .A(n486), .B(n521), .Q(\position1/N2362 ) );
  NOR21 U1043 ( .A(n487), .B(n555), .Q(\position1/N2371 ) );
  NOR21 U1044 ( .A(n487), .B(n562), .Q(\position1/N2369 ) );
  NOR21 U1045 ( .A(n487), .B(n881), .Q(\position1/N2363 ) );
  INV3 U1046 ( .A(\position1/N2352 ), .Q(n881) );
  NAND41 U1047 ( .A(n1485), .B(n1484), .C(n1483), .D(n1482), .Q(
        \position1/N2352 ) );
  NOR21 U1048 ( .A(n884), .B(n885), .Q(n1484) );
  NOR21 U1049 ( .A(n485), .B(n528), .Q(\position1/N2360 ) );
  NOR21 U1050 ( .A(n485), .B(n1100), .Q(\position1/N2354 ) );
  INV3 U1051 ( .A(\position1/N1935 ), .Q(n1100) );
  NAND41 U1052 ( .A(n1819), .B(n1818), .C(n1817), .D(n1816), .Q(
        \position1/N1935 ) );
  NOR21 U1053 ( .A(n1103), .B(n1104), .Q(n1818) );
  INV3 U1054 ( .A(n1934), .Q(n1232) );
  NAND22 U1055 ( .A(n274), .B(n1233), .Q(n1934) );
  INV3 U1056 ( .A(n1600), .Q(n1013) );
  NAND22 U1057 ( .A(n274), .B(n1014), .Q(n1600) );
  INV3 U1058 ( .A(n1936), .Q(n1236) );
  NAND22 U1059 ( .A(n628), .B(n1237), .Q(n1936) );
  INV3 U1060 ( .A(n1602), .Q(n1017) );
  NAND22 U1061 ( .A(n628), .B(n1018), .Q(n1602) );
  INV3 U1062 ( .A(\gensync1/n99 ), .Q(cam_y[0]) );
  NOR21 U1063 ( .A(n411), .B(n412), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [11]) );
  INV3 U1064 ( .A(\position1/N365 ), .Q(n412) );
  INV3 U1065 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [10]), 
        .Q(n411) );
  NOR21 U1066 ( .A(n349), .B(n412), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [11]) );
  INV3 U1067 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [10]), 
        .Q(n349) );
  NOR21 U1068 ( .A(n437), .B(n438), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [11]) );
  INV3 U1069 ( .A(\position1/N290 ), .Q(n438) );
  INV3 U1070 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [10]), 
        .Q(n437) );
  NOR21 U1071 ( .A(n365), .B(n438), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [11]) );
  INV3 U1072 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [10]), 
        .Q(n365) );
  NOR21 U1073 ( .A(n413), .B(n414), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [12]) );
  INV3 U1074 ( .A(\position1/N366 ), .Q(n414) );
  INV3 U1075 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [11]), 
        .Q(n413) );
  NOR21 U1076 ( .A(n350), .B(n414), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [12]) );
  INV3 U1077 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [11]), 
        .Q(n350) );
  NOR21 U1078 ( .A(n439), .B(n440), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [12]) );
  INV3 U1079 ( .A(\position1/N291 ), .Q(n440) );
  INV3 U1080 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [11]), 
        .Q(n439) );
  NOR21 U1081 ( .A(n366), .B(n440), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [12]) );
  INV3 U1082 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [11]), 
        .Q(n366) );
  NOR21 U1083 ( .A(n412), .B(n231), .Q(\position1/r413/carry [11]) );
  INV3 U1084 ( .A(\position1/r413/carry [10]), .Q(n231) );
  NOR21 U1085 ( .A(n416), .B(n233), .Q(\position1/r413/carry [13]) );
  INV3 U1086 ( .A(\position1/r413/carry [12]), .Q(n233) );
  NOR21 U1087 ( .A(n442), .B(n216), .Q(\position1/r412/carry [13]) );
  INV3 U1088 ( .A(\position1/r412/carry [12]), .Q(n216) );
  NOR21 U1089 ( .A(n420), .B(n235), .Q(\position1/r413/carry [15]) );
  INV3 U1090 ( .A(\position1/r413/carry [14]), .Q(n235) );
  NOR21 U1091 ( .A(n446), .B(n218), .Q(\position1/r412/carry [15]) );
  INV3 U1092 ( .A(\position1/r412/carry [14]), .Q(n218) );
  NOR21 U1093 ( .A(n424), .B(n237), .Q(\position1/r413/carry [17]) );
  INV3 U1094 ( .A(\position1/r413/carry [16]), .Q(n237) );
  NOR21 U1095 ( .A(n450), .B(n220), .Q(\position1/r412/carry [17]) );
  INV3 U1096 ( .A(\position1/r412/carry [16]), .Q(n220) );
  NOR21 U1097 ( .A(n428), .B(n239), .Q(\position1/r413/carry [19]) );
  INV3 U1098 ( .A(\position1/r413/carry [18]), .Q(n239) );
  NOR21 U1099 ( .A(n454), .B(n222), .Q(\position1/r412/carry [19]) );
  INV3 U1100 ( .A(\position1/r412/carry [18]), .Q(n222) );
  NOR21 U1101 ( .A(n432), .B(n241), .Q(\position1/r413/carry [21]) );
  INV3 U1102 ( .A(\position1/r413/carry [20]), .Q(n241) );
  NOR21 U1103 ( .A(n458), .B(n224), .Q(\position1/r412/carry [21]) );
  INV3 U1104 ( .A(\position1/r412/carry [20]), .Q(n224) );
  NOR21 U1105 ( .A(n362), .B(n243), .Q(\position1/r413/carry [23]) );
  INV3 U1106 ( .A(\position1/r413/carry [22]), .Q(n243) );
  NOR21 U1107 ( .A(n378), .B(n226), .Q(\position1/r412/carry [23]) );
  INV3 U1108 ( .A(\position1/r412/carry [22]), .Q(n226) );
  NOR21 U1109 ( .A(n414), .B(n232), .Q(\position1/r413/carry [12]) );
  INV3 U1110 ( .A(\position1/r413/carry [11]), .Q(n232) );
  NOR21 U1111 ( .A(n418), .B(n234), .Q(\position1/r413/carry [14]) );
  INV3 U1112 ( .A(\position1/r413/carry [13]), .Q(n234) );
  NOR21 U1113 ( .A(n444), .B(n217), .Q(\position1/r412/carry [14]) );
  INV3 U1114 ( .A(\position1/r412/carry [13]), .Q(n217) );
  NOR21 U1115 ( .A(n422), .B(n236), .Q(\position1/r413/carry [16]) );
  INV3 U1116 ( .A(\position1/r413/carry [15]), .Q(n236) );
  NOR21 U1117 ( .A(n448), .B(n219), .Q(\position1/r412/carry [16]) );
  INV3 U1118 ( .A(\position1/r412/carry [15]), .Q(n219) );
  NOR21 U1119 ( .A(n426), .B(n238), .Q(\position1/r413/carry [18]) );
  INV3 U1120 ( .A(\position1/r413/carry [17]), .Q(n238) );
  NOR21 U1121 ( .A(n452), .B(n221), .Q(\position1/r412/carry [18]) );
  INV3 U1122 ( .A(\position1/r412/carry [17]), .Q(n221) );
  NOR21 U1123 ( .A(n430), .B(n240), .Q(\position1/r413/carry [20]) );
  INV3 U1124 ( .A(\position1/r413/carry [19]), .Q(n240) );
  NOR21 U1125 ( .A(n456), .B(n223), .Q(\position1/r412/carry [20]) );
  INV3 U1126 ( .A(\position1/r412/carry [19]), .Q(n223) );
  NOR21 U1127 ( .A(n434), .B(n242), .Q(\position1/r413/carry [22]) );
  INV3 U1128 ( .A(\position1/r413/carry [21]), .Q(n242) );
  NOR21 U1129 ( .A(n460), .B(n225), .Q(\position1/r412/carry [22]) );
  INV3 U1130 ( .A(\position1/r412/carry [21]), .Q(n225) );
  NOR21 U1131 ( .A(n229), .B(n230), .Q(\position1/r413/carry [10]) );
  INV3 U1132 ( .A(\position1/N364 ), .Q(n229) );
  INV3 U1133 ( .A(\position1/r413/carry [9]), .Q(n230) );
  NOR21 U1134 ( .A(n212), .B(n213), .Q(\position1/r412/carry [10]) );
  INV3 U1135 ( .A(\position1/N289 ), .Q(n212) );
  INV3 U1136 ( .A(\position1/r412/carry [9]), .Q(n213) );
  BUF2 U1137 ( .A(n2134), .Q(n503) );
  BUF2 U1138 ( .A(n2134), .Q(cam_x[0]) );
  NOR21 U1139 ( .A(n228), .B(\gensync1/n99 ), .Q(\position1/r413/carry [1]) );
  INV3 U1140 ( .A(\position1/N355 ), .Q(n228) );
  NOR21 U1141 ( .A(n210), .B(n211), .Q(\position1/r412/carry [1]) );
  INV3 U1142 ( .A(n503), .Q(n211) );
  INV3 U1143 ( .A(\position1/N280 ), .Q(n210) );
  NOR21 U1144 ( .A(n211), .B(n466), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [2]) );
  INV3 U1145 ( .A(\position1/N281 ), .Q(n466) );
  NOR21 U1146 ( .A(n211), .B(n466), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [2]) );
  NOR21 U1147 ( .A(\gensync1/n99 ), .B(n467), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [2]) );
  INV3 U1148 ( .A(\position1/N356 ), .Q(n467) );
  NOR21 U1149 ( .A(\gensync1/n99 ), .B(n467), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [2]) );
  XOR21 U1150 ( .A(\position1/N379 ), .B(\position1/r413/carry [24]), .Q(
        \position1/N559 ) );
  NOR21 U1151 ( .A(n364), .B(n244), .Q(\position1/r413/carry [24]) );
  INV3 U1152 ( .A(\position1/r413/carry [23]), .Q(n244) );
  XOR21 U1153 ( .A(\position1/N304 ), .B(\position1/r412/carry [24]), .Q(
        \position1/N509 ) );
  NOR21 U1154 ( .A(n380), .B(n227), .Q(\position1/r412/carry [24]) );
  INV3 U1155 ( .A(\position1/r412/carry [23]), .Q(n227) );
  XOR21 U1156 ( .A(\position1/r412/carry [23]), .B(\position1/N303 ), .Q(
        \position1/N508 ) );
  XOR21 U1157 ( .A(\position1/N303 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [23]), .Q(
        \position1/N927 ) );
  BUF2 U1158 ( .A(n2133), .Q(n501) );
  BUF2 U1159 ( .A(n2133), .Q(cam_x[1]) );
  BUF2 U1160 ( .A(\gensync1/n100 ), .Q(n505) );
  OAI2111 U1161 ( .A(\gensync1/N72 ), .B(\gensync1/N85 ), .C(n872), .D(n869), 
        .Q(\gensync1/n100 ) );
  INV3 U1162 ( .A(\gensync1/N69 ), .Q(n869) );
  NOR21 U1163 ( .A(n417), .B(n418), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [14]) );
  INV3 U1164 ( .A(\position1/N368 ), .Q(n418) );
  INV3 U1165 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [13]), 
        .Q(n417) );
  NOR21 U1166 ( .A(n352), .B(n418), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [14]) );
  INV3 U1167 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [13]), 
        .Q(n352) );
  NOR21 U1168 ( .A(n443), .B(n444), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [14]) );
  INV3 U1169 ( .A(\position1/N293 ), .Q(n444) );
  INV3 U1170 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [13]), 
        .Q(n443) );
  NOR21 U1171 ( .A(n368), .B(n444), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [14]) );
  INV3 U1172 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [13]), 
        .Q(n368) );
  NOR21 U1173 ( .A(n421), .B(n422), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [16]) );
  INV3 U1174 ( .A(\position1/N370 ), .Q(n422) );
  INV3 U1175 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [15]), 
        .Q(n421) );
  NOR21 U1176 ( .A(n354), .B(n422), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [16]) );
  INV3 U1177 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [15]), 
        .Q(n354) );
  NOR21 U1178 ( .A(n447), .B(n448), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [16]) );
  INV3 U1179 ( .A(\position1/N295 ), .Q(n448) );
  INV3 U1180 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [15]), 
        .Q(n447) );
  NOR21 U1181 ( .A(n370), .B(n448), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [16]) );
  INV3 U1182 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [15]), 
        .Q(n370) );
  NOR21 U1183 ( .A(n425), .B(n426), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [18]) );
  INV3 U1184 ( .A(\position1/N372 ), .Q(n426) );
  INV3 U1185 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [17]), 
        .Q(n425) );
  NOR21 U1186 ( .A(n356), .B(n426), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [18]) );
  INV3 U1187 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [17]), 
        .Q(n356) );
  NOR21 U1188 ( .A(n451), .B(n452), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [18]) );
  INV3 U1189 ( .A(\position1/N297 ), .Q(n452) );
  INV3 U1190 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [17]), 
        .Q(n451) );
  NOR21 U1191 ( .A(n372), .B(n452), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [18]) );
  INV3 U1192 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [17]), 
        .Q(n372) );
  NOR21 U1193 ( .A(n429), .B(n430), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [20]) );
  INV3 U1194 ( .A(\position1/N374 ), .Q(n430) );
  INV3 U1195 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [19]), 
        .Q(n429) );
  NOR21 U1196 ( .A(n358), .B(n430), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [20]) );
  INV3 U1197 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [19]), 
        .Q(n358) );
  NOR21 U1198 ( .A(n455), .B(n456), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [20]) );
  INV3 U1199 ( .A(\position1/N299 ), .Q(n456) );
  INV3 U1200 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [19]), 
        .Q(n455) );
  NOR21 U1201 ( .A(n374), .B(n456), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [20]) );
  INV3 U1202 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [19]), 
        .Q(n374) );
  NOR21 U1203 ( .A(n433), .B(n434), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [22]) );
  INV3 U1204 ( .A(\position1/N376 ), .Q(n434) );
  INV3 U1205 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [21]), 
        .Q(n433) );
  NOR21 U1206 ( .A(n360), .B(n434), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [22]) );
  INV3 U1207 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [21]), 
        .Q(n360) );
  NOR21 U1208 ( .A(n459), .B(n460), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [22]) );
  INV3 U1209 ( .A(\position1/N301 ), .Q(n460) );
  INV3 U1210 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [21]), 
        .Q(n459) );
  NOR21 U1211 ( .A(n376), .B(n460), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [22]) );
  INV3 U1212 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [21]), 
        .Q(n376) );
  NOR21 U1213 ( .A(n436), .B(n364), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [24]) );
  INV3 U1214 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [23]), 
        .Q(n436) );
  NOR21 U1215 ( .A(n462), .B(n380), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [24]) );
  INV3 U1216 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [23]), 
        .Q(n462) );
  XOR21 U1217 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [24]), 
        .B(\position1/N379 ), .Q(\position1/N1003 ) );
  NOR21 U1218 ( .A(n363), .B(n364), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [24]) );
  INV3 U1219 ( .A(\position1/N378 ), .Q(n364) );
  INV3 U1220 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [23]), 
        .Q(n363) );
  XOR21 U1221 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [24]), 
        .B(\position1/N304 ), .Q(\position1/N928 ) );
  NOR21 U1222 ( .A(n379), .B(n380), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [24]) );
  INV3 U1223 ( .A(\position1/N303 ), .Q(n380) );
  INV3 U1224 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [23]), 
        .Q(n379) );
  NOR21 U1225 ( .A(n415), .B(n416), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [13]) );
  INV3 U1226 ( .A(\position1/N367 ), .Q(n416) );
  INV3 U1227 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [12]), 
        .Q(n415) );
  NOR21 U1228 ( .A(n351), .B(n416), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [13]) );
  INV3 U1229 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [12]), 
        .Q(n351) );
  NOR21 U1230 ( .A(n441), .B(n442), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [13]) );
  INV3 U1231 ( .A(\position1/N292 ), .Q(n442) );
  INV3 U1232 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [12]), 
        .Q(n441) );
  NOR21 U1233 ( .A(n367), .B(n442), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [13]) );
  INV3 U1234 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [12]), 
        .Q(n367) );
  NOR21 U1235 ( .A(n419), .B(n420), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [15]) );
  INV3 U1236 ( .A(\position1/N369 ), .Q(n420) );
  INV3 U1237 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [14]), 
        .Q(n419) );
  NOR21 U1238 ( .A(n353), .B(n420), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [15]) );
  INV3 U1239 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [14]), 
        .Q(n353) );
  NOR21 U1240 ( .A(n445), .B(n446), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [15]) );
  INV3 U1241 ( .A(\position1/N294 ), .Q(n446) );
  INV3 U1242 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [14]), 
        .Q(n445) );
  NOR21 U1243 ( .A(n369), .B(n446), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [15]) );
  INV3 U1244 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [14]), 
        .Q(n369) );
  NOR21 U1245 ( .A(n423), .B(n424), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [17]) );
  INV3 U1246 ( .A(\position1/N371 ), .Q(n424) );
  INV3 U1247 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [16]), 
        .Q(n423) );
  NOR21 U1248 ( .A(n355), .B(n424), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [17]) );
  INV3 U1249 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [16]), 
        .Q(n355) );
  NOR21 U1250 ( .A(n449), .B(n450), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [17]) );
  INV3 U1251 ( .A(\position1/N296 ), .Q(n450) );
  INV3 U1252 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [16]), 
        .Q(n449) );
  NOR21 U1253 ( .A(n371), .B(n450), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [17]) );
  INV3 U1254 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [16]), 
        .Q(n371) );
  NOR21 U1255 ( .A(n427), .B(n428), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [19]) );
  INV3 U1256 ( .A(\position1/N373 ), .Q(n428) );
  INV3 U1257 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [18]), 
        .Q(n427) );
  NOR21 U1258 ( .A(n357), .B(n428), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [19]) );
  INV3 U1259 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [18]), 
        .Q(n357) );
  NOR21 U1260 ( .A(n453), .B(n454), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [19]) );
  INV3 U1261 ( .A(\position1/N298 ), .Q(n454) );
  INV3 U1262 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [18]), 
        .Q(n453) );
  NOR21 U1263 ( .A(n373), .B(n454), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [19]) );
  INV3 U1264 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [18]), 
        .Q(n373) );
  NOR21 U1265 ( .A(n431), .B(n432), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [21]) );
  INV3 U1266 ( .A(\position1/N375 ), .Q(n432) );
  INV3 U1267 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [20]), 
        .Q(n431) );
  NOR21 U1268 ( .A(n359), .B(n432), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [21]) );
  INV3 U1269 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [20]), 
        .Q(n359) );
  NOR21 U1270 ( .A(n457), .B(n458), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [21]) );
  INV3 U1271 ( .A(\position1/N300 ), .Q(n458) );
  INV3 U1272 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [20]), 
        .Q(n457) );
  NOR21 U1273 ( .A(n375), .B(n458), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [21]) );
  INV3 U1274 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [20]), 
        .Q(n375) );
  NOR21 U1275 ( .A(n435), .B(n362), .Q(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [23]) );
  INV3 U1276 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [22]), 
        .Q(n435) );
  NOR21 U1277 ( .A(n361), .B(n362), .Q(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [23]) );
  INV3 U1278 ( .A(\position1/N377 ), .Q(n362) );
  INV3 U1279 ( .A(\position1/dp_cluster_2/add_0_root_add_189_3/carry [22]), 
        .Q(n361) );
  NOR21 U1280 ( .A(n461), .B(n378), .Q(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [23]) );
  INV3 U1281 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [22]), 
        .Q(n461) );
  NOR21 U1282 ( .A(n377), .B(n378), .Q(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [23]) );
  INV3 U1283 ( .A(\position1/N302 ), .Q(n378) );
  INV3 U1284 ( .A(\position1/dp_cluster_3/add_0_root_add_188_3/carry [22]), 
        .Q(n377) );
  NOR21 U1285 ( .A(n440), .B(n215), .Q(\position1/r412/carry [12]) );
  INV3 U1286 ( .A(\position1/r412/carry [11]), .Q(n215) );
  NOR21 U1287 ( .A(n438), .B(n214), .Q(\position1/r412/carry [11]) );
  INV3 U1288 ( .A(\position1/r412/carry [10]), .Q(n214) );
  BUF2 U1289 ( .A(n2132), .Q(n499) );
  XOR21 U1290 ( .A(\position1/r413/carry [23]), .B(\position1/N378 ), .Q(
        \position1/N558 ) );
  XOR21 U1291 ( .A(\position1/r413/carry [22]), .B(\position1/N377 ), .Q(
        \position1/N557 ) );
  XOR21 U1292 ( .A(\position1/r412/carry [21]), .B(\position1/N301 ), .Q(
        \position1/N506 ) );
  XOR21 U1293 ( .A(\position1/r412/carry [22]), .B(\position1/N302 ), .Q(
        \position1/N507 ) );
  XOR21 U1294 ( .A(\position1/N378 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [23]), .Q(
        \position1/N1002 ) );
  XOR21 U1295 ( .A(\position1/N376 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [21]), .Q(
        \position1/N1000 ) );
  XOR21 U1296 ( .A(\position1/N377 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [22]), .Q(
        \position1/N1001 ) );
  XOR21 U1297 ( .A(\position1/N301 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [21]), .Q(
        \position1/N925 ) );
  XOR21 U1298 ( .A(\position1/N302 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [22]), .Q(
        \position1/N926 ) );
  BUF2 U1299 ( .A(n2132), .Q(cam_x[2]) );
  BUF2 U1300 ( .A(n2131), .Q(cam_x[3]) );
  INV3 U1301 ( .A(\position1/dp_cluster_5/add_179_aco/carry [23]), .Q(n410) );
  INV3 U1302 ( .A(\position1/dp_cluster_4/add_178_aco/carry [23]), .Q(n395) );
  INV3 U1303 ( .A(\position1/n1151 ), .Q(n1361) );
  INV3 U1304 ( .A(\position1/n1145 ), .Q(n1360) );
  XOR21 U1305 ( .A(\position1/r413/carry [19]), .B(\position1/N374 ), .Q(
        \position1/N554 ) );
  XOR21 U1306 ( .A(\position1/r413/carry [20]), .B(\position1/N375 ), .Q(
        \position1/N555 ) );
  XOR21 U1307 ( .A(\position1/r413/carry [21]), .B(\position1/N376 ), .Q(
        \position1/N556 ) );
  XOR21 U1308 ( .A(\position1/r412/carry [18]), .B(\position1/N298 ), .Q(
        \position1/N503 ) );
  XOR21 U1309 ( .A(\position1/r412/carry [19]), .B(\position1/N299 ), .Q(
        \position1/N504 ) );
  XOR21 U1310 ( .A(\position1/r412/carry [20]), .B(\position1/N300 ), .Q(
        \position1/N505 ) );
  XOR21 U1311 ( .A(\position1/N374 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [19]), .Q(
        \position1/N998 ) );
  XOR21 U1312 ( .A(\position1/N375 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [20]), .Q(
        \position1/N999 ) );
  XOR21 U1313 ( .A(\position1/N298 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [18]), .Q(
        \position1/N922 ) );
  XOR21 U1314 ( .A(\position1/N299 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [19]), .Q(
        \position1/N923 ) );
  XOR21 U1315 ( .A(\position1/N300 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [20]), .Q(
        \position1/N924 ) );
  NOR21 U1316 ( .A(n505), .B(n7), .Q(n2130) );
  BUF2 U1317 ( .A(n2131), .Q(n497) );
  INV3 U1318 ( .A(\gensync1/n94 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [6]) );
  NOR21 U1319 ( .A(n505), .B(n6), .Q(n2128) );
  XOR21 U1320 ( .A(\position1/r413/carry [17]), .B(\position1/N372 ), .Q(
        \position1/N552 ) );
  XOR21 U1321 ( .A(\position1/r413/carry [18]), .B(\position1/N373 ), .Q(
        \position1/N553 ) );
  XOR21 U1322 ( .A(\position1/r412/carry [16]), .B(\position1/N296 ), .Q(
        \position1/N501 ) );
  XOR21 U1323 ( .A(\position1/r412/carry [17]), .B(\position1/N297 ), .Q(
        \position1/N502 ) );
  XOR21 U1324 ( .A(\position1/N372 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [17]), .Q(
        \position1/N996 ) );
  XOR21 U1325 ( .A(\position1/N373 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [18]), .Q(
        \position1/N997 ) );
  XOR21 U1326 ( .A(\position1/N296 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [16]), .Q(
        \position1/N920 ) );
  XOR21 U1327 ( .A(\position1/N297 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [17]), .Q(
        \position1/N921 ) );
  BUF2 U1328 ( .A(n2129), .Q(n493) );
  BUF2 U1329 ( .A(n2129), .Q(cam_x[5]) );
  XOR21 U1330 ( .A(\position1/r413/carry [14]), .B(\position1/N369 ), .Q(
        \position1/N549 ) );
  XOR21 U1331 ( .A(\position1/r413/carry [15]), .B(\position1/N370 ), .Q(
        \position1/N550 ) );
  XOR21 U1332 ( .A(\position1/r413/carry [16]), .B(\position1/N371 ), .Q(
        \position1/N551 ) );
  XOR21 U1333 ( .A(\position1/r412/carry [14]), .B(\position1/N294 ), .Q(
        \position1/N499 ) );
  XOR21 U1334 ( .A(\position1/r412/carry [15]), .B(\position1/N295 ), .Q(
        \position1/N500 ) );
  XOR21 U1335 ( .A(\position1/N370 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [15]), .Q(
        \position1/N994 ) );
  XOR21 U1336 ( .A(\position1/N371 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [16]), .Q(
        \position1/N995 ) );
  XOR21 U1337 ( .A(\position1/N294 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [14]), .Q(
        \position1/N918 ) );
  XOR21 U1338 ( .A(\position1/N295 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [15]), .Q(
        \position1/N919 ) );
  BUF2 U1339 ( .A(n2127), .Q(cam_x[7]) );
  XOR21 U1340 ( .A(\position1/r413/carry [12]), .B(\position1/N367 ), .Q(
        \position1/N547 ) );
  XOR21 U1341 ( .A(\position1/r413/carry [13]), .B(\position1/N368 ), .Q(
        \position1/N548 ) );
  XOR21 U1342 ( .A(\position1/r412/carry [11]), .B(\position1/N291 ), .Q(
        \position1/N496 ) );
  XOR21 U1343 ( .A(\position1/r412/carry [12]), .B(\position1/N292 ), .Q(
        \position1/N497 ) );
  XOR21 U1344 ( .A(\position1/r412/carry [13]), .B(\position1/N293 ), .Q(
        \position1/N498 ) );
  XOR21 U1345 ( .A(\position1/N367 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [12]), .Q(
        \position1/N991 ) );
  XOR21 U1346 ( .A(\position1/N368 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [13]), .Q(
        \position1/N992 ) );
  XOR21 U1347 ( .A(\position1/N369 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [14]), .Q(
        \position1/N993 ) );
  XOR21 U1348 ( .A(\position1/N292 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [12]), .Q(
        \position1/N916 ) );
  XOR21 U1349 ( .A(\position1/N293 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [13]), .Q(
        \position1/N917 ) );
  BUF2 U1350 ( .A(n2127), .Q(n489) );
  AOI221 U1351 ( .A(\position1/N338 ), .B(n644), .C(\position1/N615 ), .D(n645), .Q(\position1/n1020 ) );
  AOI221 U1352 ( .A(\position1/N545 ), .B(n512), .C(\position1/N989 ), .D(n640), .Q(\position1/n914 ) );
  XOR21 U1353 ( .A(\position1/N365 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [10]), .Q(
        \position1/N989 ) );
  XOR21 U1354 ( .A(\position1/r413/carry [10]), .B(\position1/N365 ), .Q(
        \position1/N545 ) );
  XOR21 U1355 ( .A(\position1/N365 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [10]), .Q(
        \position1/N415 ) );
  XOR21 U1356 ( .A(\position1/r413/carry [9]), .B(\position1/N364 ), .Q(
        \position1/N544 ) );
  XOR21 U1357 ( .A(\position1/r412/carry [9]), .B(\position1/N289 ), .Q(
        \position1/N494 ) );
  XOR21 U1358 ( .A(\position1/r413/carry [11]), .B(\position1/N366 ), .Q(
        \position1/N546 ) );
  XOR21 U1359 ( .A(\position1/r412/carry [10]), .B(\position1/N290 ), .Q(
        \position1/N495 ) );
  XOR21 U1360 ( .A(\position1/N366 ), .B(
        \position1/dp_cluster_2/add_0_root_add_189_3/carry [11]), .Q(
        \position1/N990 ) );
  XOR21 U1361 ( .A(\position1/N290 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [10]), .Q(
        \position1/N914 ) );
  XOR21 U1362 ( .A(\position1/N291 ), .B(
        \position1/dp_cluster_3/add_0_root_add_188_3/carry [11]), .Q(
        \position1/N915 ) );
  INV3 U1363 ( .A(\position1/n1073 ), .Q(n671) );
  AOI221 U1364 ( .A(n633), .B(n593), .C(\position1/n1074 ), .D(n741), .Q(
        \position1/n1073 ) );
  NAND22 U1365 ( .A(\position1/n1075 ), .B(\position1/n1076 ), .Q(
        \position1/n1074 ) );
  AOI221 U1366 ( .A(n594), .B(n477), .C(\position1/N446 ), .D(n476), .Q(
        \position1/n1076 ) );
  AOI221 U1367 ( .A(\position1/N412 ), .B(n643), .C(\position1/N639 ), .D(n647), .Q(\position1/n924 ) );
  AOI221 U1368 ( .A(\position1/N413 ), .B(n643), .C(\position1/N640 ), .D(n647), .Q(\position1/n920 ) );
  AOI221 U1369 ( .A(\position1/N337 ), .B(n644), .C(\position1/N614 ), .D(n645), .Q(\position1/n1024 ) );
  AOI221 U1370 ( .A(\position1/N605 ), .B(n479), .C(\position1/N576 ), .D(n478), .Q(\position1/n1075 ) );
  XOR21 U1371 ( .A(\position1/r458/carry [16]), .B(n592), .Q(\position1/N576 )
         );
  AOI221 U1372 ( .A(\position1/N411 ), .B(n643), .C(\position1/N638 ), .D(n645), .Q(\position1/n928 ) );
  AOI221 U1373 ( .A(\position1/N335 ), .B(n643), .C(\position1/N612 ), .D(n645), .Q(\position1/n1032 ) );
  AOI221 U1374 ( .A(\position1/N336 ), .B(n642), .C(\position1/N613 ), .D(n645), .Q(\position1/n1028 ) );
  AOI221 U1375 ( .A(\position1/N603 ), .B(n479), .C(\position1/N574 ), .D(n478), .Q(\position1/n1083 ) );
  XOR21 U1376 ( .A(\position1/r458/carry [14]), .B(n475), .Q(\position1/N574 )
         );
  AOI221 U1377 ( .A(\position1/N604 ), .B(n479), .C(\position1/N575 ), .D(n478), .Q(\position1/n1079 ) );
  XOR21 U1378 ( .A(\position1/r458/carry [15]), .B(n596), .Q(\position1/N575 )
         );
  INV3 U1379 ( .A(\position1/n1081 ), .Q(n669) );
  AOI221 U1380 ( .A(n633), .B(\position1/N2447 ), .C(\position1/n1082 ), .D(
        n741), .Q(\position1/n1081 ) );
  NAND22 U1381 ( .A(\position1/n1083 ), .B(\position1/n1084 ), .Q(
        \position1/n1082 ) );
  AOI221 U1382 ( .A(\position1/N2447 ), .B(n477), .C(\position1/N444 ), .D(
        n476), .Q(\position1/n1084 ) );
  INV3 U1383 ( .A(\position1/n1077 ), .Q(n670) );
  AOI221 U1384 ( .A(n633), .B(n597), .C(\position1/n1078 ), .D(n741), .Q(
        \position1/n1077 ) );
  NAND22 U1385 ( .A(\position1/n1079 ), .B(\position1/n1080 ), .Q(
        \position1/n1078 ) );
  AOI221 U1386 ( .A(n598), .B(n477), .C(\position1/N445 ), .D(n476), .Q(
        \position1/n1080 ) );
  NAND22 U1387 ( .A(reset_top), .B(\position1/n1182 ), .Q(\position1/n1177 )
         );
  NAND31 U1388 ( .A(\position1/n1065 ), .B(\position1/n1149 ), .C(n781), .Q(
        \position1/n1063 ) );
  INV3 U1389 ( .A(\position1/n1062 ), .Q(n781) );
  XOR21 U1390 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), 
        .B(\position1/add_250_2/carry[4] ), .Q(\position1/N2408 ) );
  XOR21 U1391 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), 
        .B(\position1/add_250_2/carry[6] ), .Q(\position1/N2410 ) );
  XOR21 U1392 ( .A(\position1/add_250_2/carry[8] ), .B(
        \position1/dp_cluster_6/N389 ), .Q(\position1/N2412 ) );
  NOR21 U1393 ( .A(n318), .B(\gensync1/n92 ), .Q(
        \position1/add_250_2/carry[8] ) );
  INV3 U1394 ( .A(\position1/add_250_2/carry[7] ), .Q(n318) );
  XOR21 U1395 ( .A(\position1/add_250/carry[8] ), .B(
        \position1/dp_cluster_7/N314 ), .Q(\position1/N2401 ) );
  NOR21 U1396 ( .A(n313), .B(n314), .Q(\position1/add_250/carry[8] ) );
  INV3 U1397 ( .A(n489), .Q(n314) );
  INV3 U1398 ( .A(\position1/add_250/carry[7] ), .Q(n313) );
  NAND22 U1399 ( .A(\position1/n1144 ), .B(\position1/n1062 ), .Q(
        \position1/n1141 ) );
  NOR21 U1400 ( .A(\position1/n1182 ), .B(n651), .Q(\position1/n1179 ) );
  XNR21 U1401 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), 
        .B(\position1/sub_250_3/carry[7] ), .Q(\position1/N2389 ) );
  XOR21 U1402 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), 
        .B(\position1/add_250_2/carry[3] ), .Q(\position1/N2407 ) );
  BUF6 U1403 ( .A(\position1/n1060 ), .Q(n478) );
  XOR21 U1404 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), 
        .B(cam_y[0]), .Q(\position1/N2383 ) );
  XOR21 U1405 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), 
        .B(\position1/add_250_2/carry[7] ), .Q(\position1/N2411 ) );
  NOR21 U1406 ( .A(\position1/n1057 ), .B(\position1/n1058 ), .Q(
        \position1/n857 ) );
  XOR21 U1407 ( .A(n151), .B(\position1/dp_cluster_7/N314 ), .Q(
        \position1/N2380 ) );
  NOR21 U1408 ( .A(\position1/sub_250/carry[7] ), .B(n489), .Q(n151) );
  XNR21 U1409 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), 
        .B(\position1/sub_250_3/carry[4] ), .Q(\position1/N2386 ) );
  XNR21 U1410 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), 
        .B(\position1/sub_250_3/carry[6] ), .Q(\position1/N2388 ) );
  BUF6 U1411 ( .A(\position1/n1070 ), .Q(n477) );
  OAI2111 U1412 ( .A(n1361), .B(\position1/n1063 ), .C(\position1/n1142 ), .D(
        \position1/n1143 ), .Q(\position1/n1070 ) );
  NAND22 U1413 ( .A(\position1/n1062 ), .B(n1349), .Q(\position1/n1143 ) );
  NAND31 U1414 ( .A(n782), .B(\position1/n1145 ), .C(n1359), .Q(
        \position1/n1142 ) );
  XNR21 U1415 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), 
        .B(\position1/add_250_2/carry[2] ), .Q(\position1/N2406 ) );
  INV3 U1416 ( .A(\position1/n1085 ), .Q(n668) );
  AOI221 U1417 ( .A(n633), .B(n601), .C(\position1/n1086 ), .D(n741), .Q(
        \position1/n1085 ) );
  NAND22 U1418 ( .A(\position1/n1087 ), .B(\position1/n1088 ), .Q(
        \position1/n1086 ) );
  AOI221 U1419 ( .A(n602), .B(n477), .C(\position1/N443 ), .D(n476), .Q(
        \position1/n1088 ) );
  AOI221 U1420 ( .A(n516), .B(n477), .C(n513), .D(n476), .Q(\position1/n1140 )
         );
  AOI221 U1421 ( .A(n632), .B(n477), .C(\position1/N431 ), .D(n476), .Q(
        \position1/n1136 ) );
  XNR21 U1422 ( .A(n515), .B(n630), .Q(\position1/N431 ) );
  AOI221 U1423 ( .A(n627), .B(n477), .C(\position1/N432 ), .D(n476), .Q(
        \position1/n1132 ) );
  XOR21 U1424 ( .A(\position1/r457/carry[2] ), .B(n625), .Q(\position1/N432 )
         );
  AOI221 U1425 ( .A(n623), .B(n477), .C(\position1/N433 ), .D(n476), .Q(
        \position1/n1128 ) );
  XOR21 U1426 ( .A(\position1/r457/carry[3] ), .B(n621), .Q(\position1/N433 )
         );
  AOI221 U1427 ( .A(\position1/N2457 ), .B(n477), .C(\position1/N434 ), .D(
        n476), .Q(\position1/n1124 ) );
  XOR21 U1428 ( .A(\position1/r457/carry[4] ), .B(\position1/N2457 ), .Q(
        \position1/N434 ) );
  AOI221 U1429 ( .A(n620), .B(n477), .C(\position1/N435 ), .D(n476), .Q(
        \position1/n1120 ) );
  XOR21 U1430 ( .A(\position1/r457/carry[5] ), .B(n618), .Q(\position1/N435 )
         );
  AOI221 U1431 ( .A(n470), .B(n477), .C(\position1/N436 ), .D(n476), .Q(
        \position1/n1116 ) );
  XOR21 U1432 ( .A(\position1/r457/carry[6] ), .B(n470), .Q(\position1/N436 )
         );
  AOI221 U1433 ( .A(n616), .B(n477), .C(\position1/N437 ), .D(n476), .Q(
        \position1/n1112 ) );
  XOR21 U1434 ( .A(\position1/r457/carry[7] ), .B(n613), .Q(\position1/N437 )
         );
  AOI221 U1435 ( .A(\position1/N2453 ), .B(n477), .C(\position1/N438 ), .D(
        n476), .Q(\position1/n1108 ) );
  XOR21 U1436 ( .A(\position1/r457/carry[8] ), .B(\position1/N2453 ), .Q(
        \position1/N438 ) );
  AOI221 U1437 ( .A(n610), .B(n477), .C(\position1/N439 ), .D(n476), .Q(
        \position1/n1104 ) );
  XOR21 U1438 ( .A(\position1/r457/carry[9] ), .B(n607), .Q(\position1/N439 )
         );
  AOI221 U1439 ( .A(n473), .B(n477), .C(\position1/N440 ), .D(n476), .Q(
        \position1/n1100 ) );
  XOR21 U1440 ( .A(\position1/r457/carry[10] ), .B(n472), .Q(\position1/N440 )
         );
  AOI221 U1441 ( .A(n606), .B(n477), .C(\position1/N441 ), .D(n476), .Q(
        \position1/n1096 ) );
  XOR21 U1442 ( .A(\position1/r457/carry[11] ), .B(n604), .Q(\position1/N441 )
         );
  AOI221 U1443 ( .A(\position1/N2449 ), .B(n477), .C(\position1/N442 ), .D(
        n476), .Q(\position1/n1092 ) );
  XOR21 U1444 ( .A(\position1/r457/carry[12] ), .B(\position1/N2449 ), .Q(
        \position1/N442 ) );
  NOR31 U1445 ( .A(\position1/n1392 ), .B(\position1/n1393 ), .C(
        \position1/n1394 ), .Q(\position1/n1391 ) );
  NAND22 U1446 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), 
        .B(\position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .Q(
        \position1/n1394 ) );
  NAND31 U1447 ( .A(cam_y[0]), .B(\gensync1/n94 ), .C(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .Q(
        \position1/n1393 ) );
  NAND41 U1448 ( .A(\position1/dp_cluster_6/N389 ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .C(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .D(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .Q(
        \position1/n1392 ) );
  NOR31 U1449 ( .A(cam_x[7]), .B(\position1/dp_cluster_7/N314 ), .C(cam_x[6]), 
        .Q(\position1/n1400 ) );
  NAND41 U1450 ( .A(cam_x[5]), .B(cam_x[6]), .C(cam_x[7]), .D(
        \position1/dp_cluster_7/N314 ), .Q(\position1/n1395 ) );
  NAND41 U1451 ( .A(cam_x[0]), .B(cam_x[1]), .C(n499), .D(cam_x[4]), .Q(
        \position1/n1396 ) );
  INV3 U1452 ( .A(\position1/n1397 ), .Q(n851) );
  AOI221 U1453 ( .A(\position1/N602 ), .B(n479), .C(\position1/N573 ), .D(n478), .Q(\position1/n1087 ) );
  XOR21 U1454 ( .A(\position1/r458/carry [13]), .B(n600), .Q(\position1/N573 )
         );
  AOI221 U1455 ( .A(\position1/N535 ), .B(n511), .C(\position1/N355 ), .D(n639), .Q(\position1/n954 ) );
  XOR21 U1456 ( .A(cam_y[0]), .B(\position1/N355 ), .Q(\position1/N535 ) );
  AOI221 U1457 ( .A(\position1/N536 ), .B(n740), .C(\position1/N980 ), .D(n640), .Q(\position1/n950 ) );
  XOR21 U1458 ( .A(\position1/N356 ), .B(cam_y[0]), .Q(\position1/N980 ) );
  AOI221 U1459 ( .A(\position1/N485 ), .B(n740), .C(\position1/N280 ), .D(n639), .Q(\position1/n1054 ) );
  XOR21 U1460 ( .A(n503), .B(\position1/N280 ), .Q(\position1/N485 ) );
  AOI221 U1461 ( .A(\position1/N486 ), .B(n740), .C(\position1/N905 ), .D(n641), .Q(\position1/n1050 ) );
  XOR21 U1462 ( .A(\position1/N281 ), .B(n503), .Q(\position1/N905 ) );
  NOR21 U1463 ( .A(\position1/N2412 ), .B(n30), .Q(n1403) );
  NOR21 U1464 ( .A(\position1/N2401 ), .B(n29), .Q(n1418) );
  NOR21 U1465 ( .A(\position1/N2377 ), .B(n22), .Q(n1442) );
  NOR21 U1466 ( .A(\position1/N2379 ), .B(n27), .Q(n1446) );
  INV3 U1467 ( .A(n152), .Q(\position1/sub_250_3/carry[4] ) );
  NOR21 U1468 ( .A(\position1/sub_250_3/carry[3] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), .Q(n152) );
  XOR21 U1469 ( .A(n156), .B(\position1/dp_cluster_6/N389 ), .Q(
        \position1/N2390 ) );
  NOR21 U1470 ( .A(\position1/sub_250_3/carry[7] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), .Q(n156) );
  INV3 U1471 ( .A(n153), .Q(\position1/sub_250_3/carry[5] ) );
  NOR21 U1472 ( .A(\position1/sub_250_3/carry[4] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), .Q(n153) );
  INV3 U1473 ( .A(n159), .Q(\position1/add_250_2/carry[2] ) );
  NOR21 U1474 ( .A(cam_y[0]), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), .Q(n159) );
  INV3 U1475 ( .A(n155), .Q(\position1/sub_250_3/carry[7] ) );
  NOR21 U1476 ( .A(\position1/sub_250_3/carry[6] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), .Q(n155) );
  INV3 U1477 ( .A(\position1/n1137 ), .Q(n655) );
  AOI221 U1478 ( .A(n633), .B(n515), .C(\position1/n1138 ), .D(n741), .Q(
        \position1/n1137 ) );
  NAND22 U1479 ( .A(\position1/n1139 ), .B(\position1/n1140 ), .Q(
        \position1/n1138 ) );
  AOI221 U1480 ( .A(n513), .B(n479), .C(n517), .D(n478), .Q(\position1/n1139 )
         );
  INV3 U1481 ( .A(\position1/n1133 ), .Q(n656) );
  AOI221 U1482 ( .A(n634), .B(n631), .C(\position1/n1134 ), .D(n741), .Q(
        \position1/n1133 ) );
  NAND22 U1483 ( .A(\position1/n1135 ), .B(\position1/n1136 ), .Q(
        \position1/n1134 ) );
  AOI221 U1484 ( .A(\position1/N590 ), .B(n479), .C(n628), .D(n478), .Q(
        \position1/n1135 ) );
  INV3 U1485 ( .A(\position1/n1129 ), .Q(n657) );
  AOI221 U1486 ( .A(n634), .B(n626), .C(\position1/n1130 ), .D(n741), .Q(
        \position1/n1129 ) );
  NAND22 U1487 ( .A(\position1/n1131 ), .B(\position1/n1132 ), .Q(
        \position1/n1130 ) );
  AOI221 U1488 ( .A(\position1/N591 ), .B(n479), .C(\position1/N562 ), .D(n478), .Q(\position1/n1131 ) );
  INV3 U1489 ( .A(\position1/n1125 ), .Q(n658) );
  AOI221 U1490 ( .A(n634), .B(n622), .C(\position1/n1126 ), .D(n741), .Q(
        \position1/n1125 ) );
  NAND22 U1491 ( .A(\position1/n1127 ), .B(\position1/n1128 ), .Q(
        \position1/n1126 ) );
  AOI221 U1492 ( .A(\position1/N592 ), .B(n479), .C(\position1/N563 ), .D(n478), .Q(\position1/n1127 ) );
  INV3 U1493 ( .A(\position1/n1121 ), .Q(n659) );
  AOI221 U1494 ( .A(n634), .B(\position1/N2457 ), .C(\position1/n1122 ), .D(
        n741), .Q(\position1/n1121 ) );
  NAND22 U1495 ( .A(\position1/n1123 ), .B(\position1/n1124 ), .Q(
        \position1/n1122 ) );
  AOI221 U1496 ( .A(\position1/N593 ), .B(n479), .C(\position1/N564 ), .D(n478), .Q(\position1/n1123 ) );
  INV3 U1497 ( .A(\position1/n1117 ), .Q(n660) );
  AOI221 U1498 ( .A(n634), .B(n619), .C(\position1/n1118 ), .D(n741), .Q(
        \position1/n1117 ) );
  NAND22 U1499 ( .A(\position1/n1119 ), .B(\position1/n1120 ), .Q(
        \position1/n1118 ) );
  AOI221 U1500 ( .A(\position1/N594 ), .B(n479), .C(\position1/N565 ), .D(n478), .Q(\position1/n1119 ) );
  INV3 U1501 ( .A(\position1/n1113 ), .Q(n661) );
  AOI221 U1502 ( .A(n634), .B(n470), .C(\position1/n1114 ), .D(n741), .Q(
        \position1/n1113 ) );
  NAND22 U1503 ( .A(\position1/n1115 ), .B(\position1/n1116 ), .Q(
        \position1/n1114 ) );
  AOI221 U1504 ( .A(\position1/N595 ), .B(n479), .C(\position1/N566 ), .D(n478), .Q(\position1/n1115 ) );
  INV3 U1505 ( .A(\position1/n1109 ), .Q(n662) );
  AOI221 U1506 ( .A(n633), .B(n615), .C(\position1/n1110 ), .D(n741), .Q(
        \position1/n1109 ) );
  NAND22 U1507 ( .A(\position1/n1111 ), .B(\position1/n1112 ), .Q(
        \position1/n1110 ) );
  AOI221 U1508 ( .A(\position1/N596 ), .B(n479), .C(\position1/N567 ), .D(n478), .Q(\position1/n1111 ) );
  INV3 U1509 ( .A(\position1/n1105 ), .Q(n663) );
  AOI221 U1510 ( .A(n633), .B(\position1/N2453 ), .C(\position1/n1106 ), .D(
        n741), .Q(\position1/n1105 ) );
  NAND22 U1511 ( .A(\position1/n1107 ), .B(\position1/n1108 ), .Q(
        \position1/n1106 ) );
  AOI221 U1512 ( .A(\position1/N597 ), .B(n479), .C(\position1/N568 ), .D(n478), .Q(\position1/n1107 ) );
  INV3 U1513 ( .A(\position1/n1101 ), .Q(n664) );
  AOI221 U1514 ( .A(n633), .B(n610), .C(\position1/n1102 ), .D(n741), .Q(
        \position1/n1101 ) );
  NAND22 U1515 ( .A(\position1/n1103 ), .B(\position1/n1104 ), .Q(
        \position1/n1102 ) );
  AOI221 U1516 ( .A(\position1/N598 ), .B(n479), .C(\position1/N569 ), .D(n478), .Q(\position1/n1103 ) );
  INV3 U1517 ( .A(\position1/n1097 ), .Q(n665) );
  AOI221 U1518 ( .A(n633), .B(n473), .C(\position1/n1098 ), .D(n741), .Q(
        \position1/n1097 ) );
  NAND22 U1519 ( .A(\position1/n1099 ), .B(\position1/n1100 ), .Q(
        \position1/n1098 ) );
  AOI221 U1520 ( .A(\position1/N599 ), .B(n479), .C(\position1/N570 ), .D(n478), .Q(\position1/n1099 ) );
  INV3 U1521 ( .A(\position1/n1093 ), .Q(n666) );
  AOI221 U1522 ( .A(n633), .B(n605), .C(\position1/n1094 ), .D(n741), .Q(
        \position1/n1093 ) );
  NAND22 U1523 ( .A(\position1/n1095 ), .B(\position1/n1096 ), .Q(
        \position1/n1094 ) );
  AOI221 U1524 ( .A(\position1/N600 ), .B(n479), .C(\position1/N571 ), .D(n478), .Q(\position1/n1095 ) );
  INV3 U1525 ( .A(\position1/n1089 ), .Q(n667) );
  AOI221 U1526 ( .A(n633), .B(\position1/N2449 ), .C(\position1/n1090 ), .D(
        n741), .Q(\position1/n1089 ) );
  NAND22 U1527 ( .A(\position1/n1091 ), .B(\position1/n1092 ), .Q(
        \position1/n1090 ) );
  AOI221 U1528 ( .A(\position1/N601 ), .B(n479), .C(\position1/N572 ), .D(n478), .Q(\position1/n1091 ) );
  INV3 U1529 ( .A(n160), .Q(\position1/add_250_2/carry[3] ) );
  NOR21 U1530 ( .A(\position1/add_250_2/carry[2] ), .B(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), .Q(n160) );
  NOR21 U1531 ( .A(\gensync1/n99 ), .B(\gensync1/n98 ), .Q(
        \position1/sub_250_3/carry[2] ) );
  NOR21 U1532 ( .A(n305), .B(\gensync1/n97 ), .Q(
        \position1/sub_250_3/carry[3] ) );
  INV3 U1533 ( .A(\position1/sub_250_3/carry[2] ), .Q(n305) );
  NOR21 U1534 ( .A(n317), .B(\gensync1/n93 ), .Q(
        \position1/add_250_2/carry[7] ) );
  INV3 U1535 ( .A(\position1/add_250_2/carry[6] ), .Q(n317) );
  NOR21 U1536 ( .A(n315), .B(\gensync1/n95 ), .Q(
        \position1/add_250_2/carry[5] ) );
  INV3 U1537 ( .A(\position1/add_250_2/carry[4] ), .Q(n315) );
  NOR21 U1538 ( .A(n160), .B(\gensync1/n96 ), .Q(
        \position1/add_250_2/carry[4] ) );
  NOR31 U1539 ( .A(\position1/n1064 ), .B(\position1/n1062 ), .C(
        \position1/n1065 ), .Q(\position1/n858 ) );
  XOR21 U1540 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), 
        .B(\position1/sub_250_3/carry[2] ), .Q(\position1/N2384 ) );
  BUF6 U1541 ( .A(\position1/n1072 ), .Q(n479) );
  INV3 U1542 ( .A(\position1/n1061 ), .Q(n673) );
  AOI311 U1543 ( .A(n741), .B(n1349), .C(\position1/n1062 ), .D(n633), .Q(
        \position1/n1061 ) );
  NOR21 U1544 ( .A(n250), .B(n251), .Q(\position1/r457/carry[6] ) );
  INV3 U1545 ( .A(n618), .Q(n250) );
  INV3 U1546 ( .A(\position1/r457/carry[5] ), .Q(n251) );
  NOR21 U1547 ( .A(n256), .B(n257), .Q(\position1/r457/carry[9] ) );
  INV3 U1548 ( .A(\position1/N2453 ), .Q(n256) );
  INV3 U1549 ( .A(\position1/r457/carry[8] ), .Q(n257) );
  NOR21 U1550 ( .A(n286), .B(n258), .Q(\position1/r457/carry[10] ) );
  INV3 U1551 ( .A(\position1/r457/carry[9] ), .Q(n258) );
  NOR21 U1552 ( .A(n269), .B(n270), .Q(\position1/r457/carry[16] ) );
  INV3 U1553 ( .A(n596), .Q(n269) );
  INV3 U1554 ( .A(\position1/r457/carry[15] ), .Q(n270) );
  NOR21 U1555 ( .A(n248), .B(n249), .Q(\position1/r457/carry[5] ) );
  INV3 U1556 ( .A(\position1/N2457 ), .Q(n248) );
  INV3 U1557 ( .A(\position1/r457/carry[4] ), .Q(n249) );
  NOR21 U1558 ( .A(n246), .B(n247), .Q(\position1/r457/carry[4] ) );
  INV3 U1559 ( .A(n621), .Q(n246) );
  INV3 U1560 ( .A(\position1/r457/carry[3] ), .Q(n247) );
  NOR21 U1561 ( .A(n245), .B(n114), .Q(\position1/r457/carry[3] ) );
  INV3 U1562 ( .A(n625), .Q(n245) );
  XOR21 U1563 ( .A(n586), .B(\position1/r457/carry[17] ), .Q(\position1/N447 )
         );
  NOR21 U1564 ( .A(n300), .B(n271), .Q(\position1/r457/carry[17] ) );
  INV3 U1565 ( .A(\position1/r457/carry[16] ), .Q(n271) );
  XOR21 U1566 ( .A(\position1/r457/carry[16] ), .B(n592), .Q(\position1/N446 )
         );
  INV3 U1567 ( .A(n114), .Q(\position1/r457/carry[2] ) );
  NOR21 U1568 ( .A(n630), .B(n515), .Q(n114) );
  NOR21 U1569 ( .A(n265), .B(n266), .Q(\position1/r457/carry[14] ) );
  INV3 U1570 ( .A(n600), .Q(n265) );
  INV3 U1571 ( .A(\position1/r457/carry[13] ), .Q(n266) );
  NOR21 U1572 ( .A(n261), .B(n262), .Q(\position1/r457/carry[12] ) );
  INV3 U1573 ( .A(n604), .Q(n261) );
  INV3 U1574 ( .A(\position1/r457/carry[11] ), .Q(n262) );
  NOR21 U1575 ( .A(n252), .B(n253), .Q(\position1/r457/carry[7] ) );
  INV3 U1576 ( .A(n470), .Q(n252) );
  INV3 U1577 ( .A(\position1/r457/carry[6] ), .Q(n253) );
  NOR21 U1578 ( .A(n263), .B(n264), .Q(\position1/r457/carry[13] ) );
  INV3 U1579 ( .A(n474), .Q(n263) );
  INV3 U1580 ( .A(\position1/r457/carry[12] ), .Q(n264) );
  NOR21 U1581 ( .A(n267), .B(n268), .Q(\position1/r457/carry[15] ) );
  INV3 U1582 ( .A(\position1/N2447 ), .Q(n267) );
  INV3 U1583 ( .A(\position1/r457/carry[14] ), .Q(n268) );
  NOR21 U1584 ( .A(n254), .B(n255), .Q(\position1/r457/carry[8] ) );
  INV3 U1585 ( .A(n613), .Q(n254) );
  INV3 U1586 ( .A(\position1/r457/carry[7] ), .Q(n255) );
  NOR21 U1587 ( .A(n259), .B(n260), .Q(\position1/r457/carry[11] ) );
  INV3 U1588 ( .A(n472), .Q(n259) );
  INV3 U1589 ( .A(\position1/r457/carry[10] ), .Q(n260) );
  NAND41 U1590 ( .A(n872), .B(\gensync1/n104 ), .C(n814), .D(\gensync1/N85 ), 
        .Q(\gensync1/n103 ) );
  NOR21 U1591 ( .A(\gensync1/N69 ), .B(\gensync1/N72 ), .Q(\gensync1/n104 ) );
  NOR21 U1592 ( .A(n272), .B(n273), .Q(\position1/r458/carry [3]) );
  INV3 U1593 ( .A(n630), .Q(n273) );
  INV3 U1594 ( .A(n625), .Q(n272) );
  NOR21 U1595 ( .A(n274), .B(n275), .Q(\position1/r458/carry [4]) );
  INV3 U1596 ( .A(n621), .Q(n274) );
  INV3 U1597 ( .A(\position1/r458/carry [3]), .Q(n275) );
  NOR21 U1598 ( .A(n276), .B(n277), .Q(\position1/r458/carry [5]) );
  INV3 U1599 ( .A(n468), .Q(n276) );
  INV3 U1600 ( .A(\position1/r458/carry [4]), .Q(n277) );
  NOR21 U1601 ( .A(n280), .B(n281), .Q(\position1/r458/carry [7]) );
  INV3 U1602 ( .A(n469), .Q(n280) );
  INV3 U1603 ( .A(\position1/r458/carry [6]), .Q(n281) );
  NOR21 U1604 ( .A(n286), .B(n287), .Q(\position1/r458/carry [10]) );
  INV3 U1605 ( .A(n607), .Q(n286) );
  INV3 U1606 ( .A(\position1/r458/carry [9]), .Q(n287) );
  NOR21 U1607 ( .A(n288), .B(n289), .Q(\position1/r458/carry [11]) );
  INV3 U1608 ( .A(n472), .Q(n288) );
  INV3 U1609 ( .A(\position1/r458/carry [10]), .Q(n289) );
  XOR21 U1610 ( .A(\position1/N356 ), .B(cam_y[0]), .Q(\position1/N406 ) );
  XOR21 U1611 ( .A(\position1/N281 ), .B(n503), .Q(\position1/N331 ) );
  XOR21 U1612 ( .A(\position1/r457/carry[14] ), .B(\position1/N2447 ), .Q(
        \position1/N444 ) );
  XOR21 U1613 ( .A(\position1/r457/carry[15] ), .B(n596), .Q(\position1/N445 )
         );
  NOR21 U1614 ( .A(n294), .B(n295), .Q(\position1/r458/carry [14]) );
  INV3 U1615 ( .A(n600), .Q(n294) );
  INV3 U1616 ( .A(\position1/r458/carry [13]), .Q(n295) );
  NOR21 U1617 ( .A(n298), .B(n299), .Q(\position1/r458/carry [16]) );
  INV3 U1618 ( .A(n596), .Q(n298) );
  INV3 U1619 ( .A(\position1/r458/carry [15]), .Q(n299) );
  NOR21 U1620 ( .A(n278), .B(n279), .Q(\position1/r458/carry [6]) );
  INV3 U1621 ( .A(n618), .Q(n278) );
  INV3 U1622 ( .A(\position1/r458/carry [5]), .Q(n279) );
  NOR21 U1623 ( .A(n290), .B(n291), .Q(\position1/r458/carry [12]) );
  INV3 U1624 ( .A(n604), .Q(n290) );
  INV3 U1625 ( .A(\position1/r458/carry [11]), .Q(n291) );
  NOR21 U1626 ( .A(n282), .B(n283), .Q(\position1/r458/carry [8]) );
  INV3 U1627 ( .A(n613), .Q(n282) );
  INV3 U1628 ( .A(\position1/r458/carry [7]), .Q(n283) );
  NOR21 U1629 ( .A(n292), .B(n293), .Q(\position1/r458/carry [13]) );
  INV3 U1630 ( .A(n474), .Q(n292) );
  INV3 U1631 ( .A(\position1/r458/carry [12]), .Q(n293) );
  NOR21 U1632 ( .A(n296), .B(n297), .Q(\position1/r458/carry [15]) );
  INV3 U1633 ( .A(n475), .Q(n296) );
  INV3 U1634 ( .A(\position1/r458/carry [14]), .Q(n297) );
  NOR21 U1635 ( .A(n284), .B(n285), .Q(\position1/r458/carry [9]) );
  INV3 U1636 ( .A(n471), .Q(n284) );
  INV3 U1637 ( .A(\position1/r458/carry [8]), .Q(n285) );
  NOR21 U1638 ( .A(\image_process1/n117 ), .B(\gensync1/n103 ), .Q(
        \image_process1/n57 ) );
  XOR21 U1639 ( .A(\position1/r457/carry[13] ), .B(n600), .Q(\position1/N443 )
         );
  NOR41 U1640 ( .A(n775), .B(\image_process1/N59 ), .C(\image_process1/N62 ), 
        .D(\image_process1/N64 ), .Q(\image_process1/n89 ) );
  INV3 U1641 ( .A(\image_process1/n57 ), .Q(n775) );
  NOR21 U1642 ( .A(\gensync1/n103 ), .B(n774), .Q(\image_process1/n58 ) );
  INV3 U1643 ( .A(\image_process1/n117 ), .Q(n774) );
  NAND22 U1644 ( .A(\gensync1/n103 ), .B(\position1/n1176 ), .Q(
        \position1/n1175 ) );
  NOR21 U1645 ( .A(\image_process1/n97 ), .B(\image_process1/N62 ), .Q(
        \image_process1/n95 ) );
  XOR21 U1646 ( .A(\position1/r458/carry [11]), .B(n604), .Q(\position1/N571 )
         );
  XOR21 U1647 ( .A(\position1/r458/carry [12]), .B(n474), .Q(\position1/N572 )
         );
  NOR21 U1648 ( .A(\gensync1/n102 ), .B(n826), .Q(\gensync1/N30 ) );
  INV3 U1649 ( .A(\gensync1/N20 ), .Q(n826) );
  INV3 U1650 ( .A(n488), .Q(n813) );
  BUF2 U1651 ( .A(n482), .Q(n483) );
  AOI211 U1652 ( .A(n487), .B(\position1/n1175 ), .C(n653), .Q(n482) );
  NOR21 U1653 ( .A(n507), .B(n818), .Q(\gensync1/N63 ) );
  INV3 U1654 ( .A(\gensync1/N53 ), .Q(n818) );
  NOR21 U1655 ( .A(n507), .B(n817), .Q(\gensync1/N64 ) );
  INV3 U1656 ( .A(\gensync1/N54 ), .Q(n817) );
  XOR21 U1657 ( .A(\position1/r458/carry [8]), .B(n471), .Q(\position1/N568 )
         );
  XOR21 U1658 ( .A(\position1/r458/carry [9]), .B(n607), .Q(\position1/N569 )
         );
  XOR21 U1659 ( .A(\position1/r458/carry [10]), .B(n472), .Q(\position1/N570 )
         );
  INV3 U1660 ( .A(\position1/n1144 ), .Q(n1349) );
  NOR21 U1661 ( .A(\gensync1/n102 ), .B(n827), .Q(\gensync1/N29 ) );
  INV3 U1662 ( .A(\gensync1/N19 ), .Q(n827) );
  NOR21 U1663 ( .A(\gensync1/n102 ), .B(n828), .Q(\gensync1/N28 ) );
  INV3 U1664 ( .A(\gensync1/N18 ), .Q(n828) );
  NOR21 U1665 ( .A(n507), .B(n819), .Q(\gensync1/N62 ) );
  INV3 U1666 ( .A(\gensync1/N52 ), .Q(n819) );
  NOR21 U1667 ( .A(n507), .B(n820), .Q(\gensync1/N61 ) );
  INV3 U1668 ( .A(\gensync1/N51 ), .Q(n820) );
  NAND22 U1669 ( .A(\position1/n1176 ), .B(n648), .Q(\position1/n1064 ) );
  INV3 U1670 ( .A(n654), .Q(n648) );
  NAND22 U1671 ( .A(\position1/n1058 ), .B(\position1/n1146 ), .Q(
        \position1/n1056 ) );
  NOR21 U1672 ( .A(n650), .B(n486), .Q(\position1/n834 ) );
  XOR21 U1673 ( .A(\position1/r458/carry [6]), .B(n469), .Q(\position1/N566 )
         );
  XOR21 U1674 ( .A(\position1/r458/carry [7]), .B(n613), .Q(\position1/N567 )
         );
  NOR21 U1675 ( .A(\gensync1/n102 ), .B(n829), .Q(\gensync1/N27 ) );
  INV3 U1676 ( .A(\gensync1/N17 ), .Q(n829) );
  BUF2 U1677 ( .A(\position1/n1152 ), .Q(n486) );
  NOR21 U1678 ( .A(n506), .B(n821), .Q(\gensync1/N60 ) );
  INV3 U1679 ( .A(\gensync1/N50 ), .Q(n821) );
  NOR21 U1680 ( .A(\image_process1/n113 ), .B(\image_process1/N59 ), .Q(
        \image_process1/n112 ) );
  INV3 U1681 ( .A(\image_process1/N59 ), .Q(n876) );
  XOR21 U1682 ( .A(\position1/r458/carry [3]), .B(n621), .Q(\position1/N563 )
         );
  XOR21 U1683 ( .A(\position1/r458/carry [4]), .B(n468), .Q(\position1/N564 )
         );
  XOR21 U1684 ( .A(\position1/r458/carry [5]), .B(n618), .Q(\position1/N565 )
         );
  BUF2 U1685 ( .A(\position1/n1152 ), .Q(n487) );
  NOR21 U1686 ( .A(\gensync1/n102 ), .B(n830), .Q(\gensync1/N26 ) );
  INV3 U1687 ( .A(\gensync1/N16 ), .Q(n830) );
  NOR21 U1688 ( .A(\gensync1/n102 ), .B(n831), .Q(\gensync1/N25 ) );
  INV3 U1689 ( .A(\gensync1/N15 ), .Q(n831) );
  BUF2 U1690 ( .A(n101), .Q(n587) );
  NOR21 U1691 ( .A(n875), .B(\image_process1/N62 ), .Q(\image_process1/n113 )
         );
  INV3 U1692 ( .A(\image_process1/N64 ), .Q(n875) );
  BUF2 U1693 ( .A(\gensync1/n101 ), .Q(n507) );
  BUF2 U1694 ( .A(\gensync1/n101 ), .Q(n506) );
  INV3 U1695 ( .A(\gensync1/N129 ), .Q(n815) );
  NOR21 U1696 ( .A(n506), .B(n822), .Q(\gensync1/N59 ) );
  INV3 U1697 ( .A(\gensync1/N49 ), .Q(n822) );
  NOR21 U1698 ( .A(n506), .B(n823), .Q(\gensync1/N58 ) );
  INV3 U1699 ( .A(\gensync1/N48 ), .Q(n823) );
  NOR21 U1700 ( .A(n506), .B(n824), .Q(\gensync1/N57 ) );
  INV3 U1701 ( .A(\gensync1/N47 ), .Q(n824) );
  INV3 U1702 ( .A(n652), .Q(n649) );
  XOR21 U1703 ( .A(n630), .B(n625), .Q(\position1/N562 ) );
  NOR21 U1704 ( .A(\gensync1/n102 ), .B(n832), .Q(\gensync1/N24 ) );
  INV3 U1705 ( .A(\gensync1/N14 ), .Q(n832) );
  NOR21 U1706 ( .A(\gensync1/n102 ), .B(n833), .Q(\gensync1/N23 ) );
  INV3 U1707 ( .A(\gensync1/N13 ), .Q(n833) );
  INV3 U1708 ( .A(n629), .Q(n628) );
  INV3 U1709 ( .A(n514), .Q(n513) );
  INV3 U1710 ( .A(n592), .Q(n300) );
  INV3 U1711 ( .A(\position1/N1570 ), .Q(n1300) );
  AOI221 U1712 ( .A(\position1/N1569 ), .B(n44), .C(n2079), .D(n2078), .Q(
        n2080) );
  NAND22 U1713 ( .A(n593), .B(n1301), .Q(n2078) );
  INV3 U1714 ( .A(\position1/N1987 ), .Q(n1081) );
  AOI221 U1715 ( .A(\position1/N1986 ), .B(n300), .C(n1745), .D(n1744), .Q(
        n1746) );
  NAND22 U1716 ( .A(n593), .B(n1082), .Q(n1744) );
  NAND22 U1717 ( .A(\position1/N1530 ), .B(n519), .Q(\position1/n1569 ) );
  NAND22 U1718 ( .A(\position1/N1947 ), .B(n553), .Q(\position1/n1373 ) );
  NAND22 U1719 ( .A(\position1/N1532 ), .B(n519), .Q(\position1/n1567 ) );
  NAND22 U1720 ( .A(\position1/N1949 ), .B(n553), .Q(\position1/n1371 ) );
  NAND22 U1721 ( .A(\position1/N1534 ), .B(n518), .Q(\position1/n1565 ) );
  NAND22 U1722 ( .A(\position1/N1951 ), .B(n552), .Q(\position1/n1369 ) );
  NAND22 U1723 ( .A(\position1/N1536 ), .B(n518), .Q(\position1/n1563 ) );
  NAND22 U1724 ( .A(\position1/N1953 ), .B(n552), .Q(\position1/n1367 ) );
  NAND22 U1725 ( .A(\position1/N1538 ), .B(n518), .Q(\position1/n1561 ) );
  NAND22 U1726 ( .A(\position1/N1955 ), .B(n552), .Q(\position1/n1365 ) );
  NAND22 U1727 ( .A(\position1/N1540 ), .B(n518), .Q(\position1/n1559 ) );
  NAND22 U1728 ( .A(\position1/N1957 ), .B(n552), .Q(\position1/n1363 ) );
  NAND22 U1729 ( .A(\position1/N1542 ), .B(n518), .Q(\position1/n1557 ) );
  NAND22 U1730 ( .A(\position1/N1959 ), .B(n552), .Q(\position1/n1361 ) );
  NAND22 U1731 ( .A(\position1/N1544 ), .B(n518), .Q(\position1/n1555 ) );
  NAND22 U1732 ( .A(\position1/N1961 ), .B(n552), .Q(\position1/n1359 ) );
  AOI221 U1733 ( .A(n524), .B(\position1/N1581 ), .C(n522), .D(
        \position1/N1554 ), .Q(\position1/n1545 ) );
  AOI221 U1734 ( .A(n558), .B(\position1/N1998 ), .C(n556), .D(
        \position1/N1971 ), .Q(\position1/n1349 ) );
  AOI221 U1735 ( .A(n524), .B(\position1/N1580 ), .C(n522), .D(
        \position1/N1553 ), .Q(\position1/n1546 ) );
  XNR21 U1736 ( .A(\position1/N1553 ), .B(n513), .Q(\position1/N1580 ) );
  AOI221 U1737 ( .A(n558), .B(\position1/N1997 ), .C(n556), .D(
        \position1/N1970 ), .Q(\position1/n1350 ) );
  XNR21 U1738 ( .A(\position1/N1970 ), .B(n513), .Q(\position1/N1997 ) );
  AOI221 U1739 ( .A(n524), .B(\position1/N1585 ), .C(n522), .D(
        \position1/N1558 ), .Q(\position1/n1541 ) );
  AOI221 U1740 ( .A(n558), .B(\position1/N2002 ), .C(n556), .D(
        \position1/N1975 ), .Q(\position1/n1345 ) );
  AOI221 U1741 ( .A(n524), .B(\position1/N1587 ), .C(n522), .D(
        \position1/N1560 ), .Q(\position1/n1539 ) );
  AOI221 U1742 ( .A(n558), .B(\position1/N2004 ), .C(n556), .D(
        \position1/N1977 ), .Q(\position1/n1343 ) );
  AOI221 U1743 ( .A(n525), .B(\position1/N1589 ), .C(n522), .D(
        \position1/N1562 ), .Q(\position1/n1537 ) );
  AOI221 U1744 ( .A(n559), .B(\position1/N2006 ), .C(n556), .D(
        \position1/N1979 ), .Q(\position1/n1341 ) );
  AOI221 U1745 ( .A(n525), .B(\position1/N1591 ), .C(n522), .D(
        \position1/N1564 ), .Q(\position1/n1535 ) );
  AOI221 U1746 ( .A(n559), .B(\position1/N2008 ), .C(n556), .D(
        \position1/N1981 ), .Q(\position1/n1339 ) );
  AOI221 U1747 ( .A(n525), .B(\position1/N1593 ), .C(n522), .D(
        \position1/N1566 ), .Q(\position1/n1533 ) );
  AOI221 U1748 ( .A(n559), .B(\position1/N2010 ), .C(n556), .D(
        \position1/N1983 ), .Q(\position1/n1337 ) );
  AOI221 U1749 ( .A(n525), .B(\position1/N1595 ), .C(n522), .D(
        \position1/N1568 ), .Q(\position1/n1531 ) );
  AOI221 U1750 ( .A(n559), .B(\position1/N2012 ), .C(n556), .D(
        \position1/N1985 ), .Q(\position1/n1335 ) );
  AOI221 U1751 ( .A(n525), .B(\position1/N1597 ), .C(n522), .D(
        \position1/N1570 ), .Q(\position1/n1529 ) );
  AOI221 U1752 ( .A(n559), .B(\position1/N2014 ), .C(n556), .D(
        \position1/N1987 ), .Q(\position1/n1333 ) );
  AOI221 U1753 ( .A(n524), .B(\position1/N1552 ), .C(n522), .D(
        \position1/N1552 ), .Q(\position1/n1547 ) );
  AOI221 U1754 ( .A(n558), .B(\position1/N1969 ), .C(n556), .D(
        \position1/N1969 ), .Q(\position1/n1351 ) );
  AOI221 U1755 ( .A(n524), .B(\position1/N1550 ), .C(n522), .D(
        \position1/N1550 ), .Q(\position1/n1549 ) );
  AOI221 U1756 ( .A(n523), .B(\position1/N1549 ), .C(n522), .D(
        \position1/N1549 ), .Q(\position1/n1550 ) );
  AOI221 U1757 ( .A(n558), .B(\position1/N1967 ), .C(n556), .D(
        \position1/N1967 ), .Q(\position1/n1353 ) );
  AOI221 U1758 ( .A(n557), .B(\position1/N1966 ), .C(n556), .D(
        \position1/N1966 ), .Q(\position1/n1354 ) );
  AOI221 U1759 ( .A(n524), .B(\position1/N1551 ), .C(n522), .D(
        \position1/N1551 ), .Q(\position1/n1548 ) );
  AOI221 U1760 ( .A(n558), .B(\position1/N1968 ), .C(n556), .D(
        \position1/N1968 ), .Q(\position1/n1352 ) );
  AOI221 U1761 ( .A(n523), .B(\position1/N1547 ), .C(n522), .D(
        \position1/N1547 ), .Q(\position1/n1552 ) );
  AOI221 U1762 ( .A(n523), .B(\position1/N1548 ), .C(n522), .D(
        \position1/N1548 ), .Q(\position1/n1551 ) );
  AOI221 U1763 ( .A(n523), .B(\position1/N1573 ), .C(n522), .D(
        \position1/N1573 ), .Q(\position1/n1553 ) );
  AOI221 U1764 ( .A(n557), .B(\position1/N1964 ), .C(n556), .D(
        \position1/N1964 ), .Q(\position1/n1356 ) );
  AOI221 U1765 ( .A(n557), .B(\position1/N1965 ), .C(n556), .D(
        \position1/N1965 ), .Q(\position1/n1355 ) );
  AOI221 U1766 ( .A(n557), .B(\position1/N1990 ), .C(n556), .D(
        \position1/N1990 ), .Q(\position1/n1357 ) );
  INV3 U1767 ( .A(\position1/N1671 ), .Q(n1247) );
  NOR21 U1768 ( .A(\position1/N1671 ), .B(n44), .Q(n2004) );
  INV3 U1769 ( .A(\position1/N2088 ), .Q(n1028) );
  NOR21 U1770 ( .A(\position1/N2088 ), .B(n300), .Q(n1670) );
  AOI221 U1771 ( .A(n524), .B(\position1/N1583 ), .C(n522), .D(
        \position1/N1556 ), .Q(\position1/n1543 ) );
  AOI221 U1772 ( .A(n558), .B(\position1/N2000 ), .C(n556), .D(
        \position1/N1973 ), .Q(\position1/n1347 ) );
  AOI221 U1773 ( .A(n1190), .B(n1928), .C(n44), .D(n1191), .Q(n1932) );
  INV3 U1774 ( .A(n1895), .Q(n1190) );
  AOI221 U1775 ( .A(\position1/n1485 ), .B(n597), .C(n1184), .D(n1193), .Q(
        n1928) );
  NOR21 U1776 ( .A(n1191), .B(n300), .Q(n1895) );
  AOI221 U1777 ( .A(n971), .B(n1594), .C(n44), .D(n972), .Q(n1598) );
  INV3 U1778 ( .A(n1561), .Q(n971) );
  AOI221 U1779 ( .A(\position1/n1289 ), .B(n597), .C(n965), .D(n974), .Q(n1594) );
  NOR21 U1780 ( .A(n972), .B(n300), .Q(n1561) );
  OAI2111 U1781 ( .A(\position1/n1436 ), .B(n594), .C(n1852), .D(n1851), .Q(
        n1853) );
  NAND22 U1782 ( .A(n298), .B(n1134), .Q(n1852) );
  OAI2111 U1783 ( .A(n296), .B(n1135), .C(n1124), .D(n1850), .Q(n1851) );
  INV3 U1784 ( .A(n1821), .Q(n1124) );
  OAI2111 U1785 ( .A(\position1/n1240 ), .B(n594), .C(n1518), .D(n1517), .Q(
        n1519) );
  NAND22 U1786 ( .A(n269), .B(n915), .Q(n1518) );
  OAI2111 U1787 ( .A(n267), .B(n916), .C(n905), .D(n1516), .Q(n1517) );
  INV3 U1788 ( .A(n1487), .Q(n905) );
  OAI2111 U1789 ( .A(\position1/n1254 ), .B(n627), .C(n1495), .D(n1494), .Q(
        n1496) );
  NAND22 U1790 ( .A(n273), .B(n936), .Q(n1495) );
  OAI2111 U1791 ( .A(n34), .B(n939), .C(n935), .D(n937), .Q(n1494) );
  INV3 U1792 ( .A(n1492), .Q(n935) );
  OAI2111 U1793 ( .A(\position1/n1252 ), .B(\position1/N2457 ), .C(n1498), .D(
        n1497), .Q(n1499) );
  NAND22 U1794 ( .A(n246), .B(n933), .Q(n1498) );
  OAI2111 U1795 ( .A(n66), .B(n934), .C(n932), .D(n1496), .Q(n1497) );
  INV3 U1796 ( .A(n1491), .Q(n932) );
  OAI2111 U1797 ( .A(\position1/n1250 ), .B(n470), .C(n1501), .D(n1500), .Q(
        n1502) );
  NAND22 U1798 ( .A(n278), .B(n930), .Q(n1501) );
  OAI2111 U1799 ( .A(n248), .B(n931), .C(n929), .D(n1499), .Q(n1500) );
  INV3 U1800 ( .A(n1490), .Q(n929) );
  OAI2111 U1801 ( .A(\position1/n1440 ), .B(n474), .C(n1846), .D(n1845), .Q(
        n1847) );
  NAND22 U1802 ( .A(n261), .B(n1140), .Q(n1846) );
  OAI2111 U1803 ( .A(n259), .B(n1142), .C(n1139), .D(n1141), .Q(n1845) );
  INV3 U1804 ( .A(n1823), .Q(n1139) );
  OAI2111 U1805 ( .A(\position1/n1244 ), .B(\position1/N2449 ), .C(n1512), .D(
        n1511), .Q(n1513) );
  NAND22 U1806 ( .A(n290), .B(n921), .Q(n1512) );
  OAI2111 U1807 ( .A(n259), .B(n923), .C(n920), .D(n922), .Q(n1511) );
  INV3 U1808 ( .A(n1489), .Q(n920) );
  OAI2111 U1809 ( .A(\position1/n1446 ), .B(n469), .C(n1835), .D(n1834), .Q(
        n1836) );
  NAND22 U1810 ( .A(n250), .B(n1149), .Q(n1835) );
  OAI2111 U1811 ( .A(n276), .B(n1150), .C(n1148), .D(n1833), .Q(n1834) );
  INV3 U1812 ( .A(n1824), .Q(n1148) );
  OAI2111 U1813 ( .A(\position1/n1438 ), .B(n475), .C(n1849), .D(n1848), .Q(
        n1850) );
  NAND22 U1814 ( .A(n294), .B(n1137), .Q(n1849) );
  OAI2111 U1815 ( .A(n292), .B(n1138), .C(n1136), .D(n1847), .Q(n1848) );
  INV3 U1816 ( .A(n1822), .Q(n1136) );
  OAI2111 U1817 ( .A(\position1/n1242 ), .B(\position1/N2447 ), .C(n1515), .D(
        n1514), .Q(n1516) );
  NAND22 U1818 ( .A(n265), .B(n918), .Q(n1515) );
  OAI2111 U1819 ( .A(n263), .B(n919), .C(n917), .D(n1513), .Q(n1514) );
  INV3 U1820 ( .A(n1488), .Q(n917) );
  OAI2111 U1821 ( .A(\position1/n1448 ), .B(n468), .C(n1832), .D(n1831), .Q(
        n1833) );
  NAND22 U1822 ( .A(n274), .B(n1152), .Q(n1832) );
  OAI2111 U1823 ( .A(n66), .B(n1153), .C(n1151), .D(n1830), .Q(n1831) );
  INV3 U1824 ( .A(n1825), .Q(n1151) );
  OAI2111 U1825 ( .A(\position1/n1450 ), .B(n627), .C(n1829), .D(n1828), .Q(
        n1830) );
  NAND22 U1826 ( .A(n273), .B(n1155), .Q(n1829) );
  OAI2111 U1827 ( .A(n513), .B(n1158), .C(n1154), .D(n1156), .Q(n1828) );
  INV3 U1828 ( .A(n1826), .Q(n1154) );
  INV3 U1829 ( .A(n1937), .Q(n1238) );
  NOR40 U1830 ( .A(n1240), .B(n1241), .C(n1242), .D(n1243), .Q(n1938) );
  NAND22 U1831 ( .A(\position1/n1524 ), .B(n515), .Q(n1937) );
  INV3 U1832 ( .A(n1603), .Q(n1019) );
  NOR40 U1833 ( .A(n1021), .B(n1022), .C(n1023), .D(n1024), .Q(n1604) );
  NAND22 U1834 ( .A(\position1/n1328 ), .B(n515), .Q(n1603) );
  NOR21 U1835 ( .A(n622), .B(\position1/n1544 ), .Q(n2016) );
  INV3 U1836 ( .A(n2008), .Q(n1295) );
  NOR21 U1837 ( .A(n621), .B(\position1/n1348 ), .Q(n1682) );
  INV3 U1838 ( .A(n1674), .Q(n1076) );
  INV3 U1839 ( .A(n1935), .Q(n1234) );
  NAND22 U1840 ( .A(\position1/n1522 ), .B(n625), .Q(n1935) );
  INV3 U1841 ( .A(n1601), .Q(n1015) );
  NAND22 U1842 ( .A(\position1/n1326 ), .B(n625), .Q(n1601) );
  INV3 U1843 ( .A(n1933), .Q(n1230) );
  NAND22 U1844 ( .A(\position1/n1520 ), .B(n468), .Q(n1933) );
  INV3 U1845 ( .A(n1599), .Q(n1011) );
  NAND22 U1846 ( .A(\position1/n1324 ), .B(\position1/N2457 ), .Q(n1599) );
  AOI2111 U1847 ( .A(n593), .B(\position1/n1436 ), .C(n1131), .D(n1123), .Q(
        n1855) );
  INV3 U1848 ( .A(n1820), .Q(n1131) );
  INV3 U1849 ( .A(n1853), .Q(n1123) );
  NAND22 U1850 ( .A(\position1/n1435 ), .B(n586), .Q(n1820) );
  AOI2111 U1851 ( .A(n591), .B(\position1/n1240 ), .C(n912), .D(n904), .Q(
        n1521) );
  INV3 U1852 ( .A(n1486), .Q(n912) );
  INV3 U1853 ( .A(n1519), .Q(n904) );
  NAND22 U1854 ( .A(\position1/n1239 ), .B(n586), .Q(n1486) );
  AOI221 U1855 ( .A(n1966), .B(n1965), .C(n44), .D(n1217), .Q(n1969) );
  NAND22 U1856 ( .A(\position1/n1508 ), .B(n592), .Q(n1966) );
  AOI221 U1857 ( .A(\position1/n1509 ), .B(n597), .C(n1964), .D(n1963), .Q(
        n1965) );
  NAND22 U1858 ( .A(n67), .B(n1218), .Q(n1964) );
  AOI221 U1859 ( .A(n1632), .B(n1631), .C(n44), .D(n998), .Q(n1635) );
  NAND22 U1860 ( .A(\position1/n1312 ), .B(n592), .Q(n1632) );
  AOI221 U1861 ( .A(\position1/n1313 ), .B(n595), .C(n1630), .D(n1629), .Q(
        n1631) );
  NAND22 U1862 ( .A(n298), .B(n999), .Q(n1630) );
  NOR21 U1863 ( .A(n1208), .B(n34), .Q(n1897) );
  NOR31 U1864 ( .A(n1211), .B(n1209), .C(n1210), .Q(n1898) );
  NOR21 U1865 ( .A(n989), .B(n34), .Q(n1563) );
  NOR31 U1866 ( .A(n992), .B(n990), .C(n991), .Q(n1564) );
  NOR21 U1867 ( .A(n1206), .B(n272), .Q(n1902) );
  NOR21 U1868 ( .A(n630), .B(\position1/n1499 ), .Q(n1900) );
  NOR21 U1869 ( .A(n987), .B(n245), .Q(n1568) );
  NOR21 U1870 ( .A(n630), .B(\position1/n1303 ), .Q(n1566) );
  NOR21 U1871 ( .A(n1204), .B(n276), .Q(n1906) );
  NOR21 U1872 ( .A(n621), .B(\position1/n1497 ), .Q(n1904) );
  NOR21 U1873 ( .A(n985), .B(n41), .Q(n1572) );
  NOR21 U1874 ( .A(n621), .B(\position1/n1301 ), .Q(n1570) );
  NOR21 U1875 ( .A(n1202), .B(n45), .Q(n1910) );
  NOR21 U1876 ( .A(n619), .B(\position1/n1495 ), .Q(n1908) );
  NOR21 U1877 ( .A(n983), .B(n252), .Q(n1576) );
  NOR21 U1878 ( .A(n618), .B(\position1/n1299 ), .Q(n1574) );
  NOR21 U1879 ( .A(n1200), .B(n284), .Q(n1914) );
  NOR21 U1880 ( .A(n614), .B(\position1/n1493 ), .Q(n1912) );
  NOR21 U1881 ( .A(n981), .B(n40), .Q(n1580) );
  NOR21 U1882 ( .A(n613), .B(\position1/n1297 ), .Q(n1578) );
  NOR21 U1883 ( .A(n1198), .B(n46), .Q(n1918) );
  NOR21 U1884 ( .A(n608), .B(\position1/n1491 ), .Q(n1916) );
  NOR21 U1885 ( .A(n979), .B(n288), .Q(n1584) );
  NOR21 U1886 ( .A(n608), .B(\position1/n1295 ), .Q(n1582) );
  AOI221 U1887 ( .A(\position1/n1542 ), .B(n620), .C(n2020), .D(n2019), .Q(
        n2021) );
  NAND22 U1888 ( .A(n278), .B(n1288), .Q(n2020) );
  AOI221 U1889 ( .A(n2018), .B(n1290), .C(n248), .D(n1291), .Q(n2019) );
  INV3 U1890 ( .A(n2017), .Q(n1290) );
  AOI221 U1891 ( .A(\position1/n1346 ), .B(n617), .C(n1686), .D(n1685), .Q(
        n1687) );
  NAND22 U1892 ( .A(n250), .B(n1069), .Q(n1686) );
  AOI221 U1893 ( .A(n1684), .B(n1071), .C(n248), .D(n1072), .Q(n1685) );
  INV3 U1894 ( .A(n1683), .Q(n1071) );
  AOI221 U1895 ( .A(\position1/n1540 ), .B(n615), .C(n2024), .D(n2023), .Q(
        n2025) );
  NAND22 U1896 ( .A(n282), .B(n1284), .Q(n2024) );
  AOI221 U1897 ( .A(n2022), .B(n2021), .C(n280), .D(n1286), .Q(n2023) );
  NAND22 U1898 ( .A(\position1/n1541 ), .B(n469), .Q(n2022) );
  AOI221 U1899 ( .A(\position1/n1344 ), .B(n615), .C(n1690), .D(n1689), .Q(
        n1691) );
  NAND22 U1900 ( .A(n254), .B(n1065), .Q(n1690) );
  AOI221 U1901 ( .A(n1688), .B(n1687), .C(n252), .D(n1067), .Q(n1689) );
  NAND22 U1902 ( .A(\position1/n1345 ), .B(n470), .Q(n1688) );
  AOI221 U1903 ( .A(\position1/n1538 ), .B(n610), .C(n2028), .D(n2027), .Q(
        n2029) );
  NAND22 U1904 ( .A(n286), .B(n1280), .Q(n2028) );
  AOI221 U1905 ( .A(n2026), .B(n2025), .C(n284), .D(n1282), .Q(n2027) );
  NAND22 U1906 ( .A(\position1/n1539 ), .B(n471), .Q(n2026) );
  AOI221 U1907 ( .A(\position1/n1342 ), .B(n609), .C(n1694), .D(n1693), .Q(
        n1695) );
  NAND22 U1908 ( .A(n286), .B(n1061), .Q(n1694) );
  AOI221 U1909 ( .A(n1692), .B(n1691), .C(n256), .D(n1063), .Q(n1693) );
  NAND22 U1910 ( .A(\position1/n1343 ), .B(n471), .Q(n1692) );
  AOI221 U1911 ( .A(\position1/n1536 ), .B(n605), .C(n2032), .D(n2031), .Q(
        n2033) );
  NAND22 U1912 ( .A(n38), .B(n1276), .Q(n2032) );
  AOI221 U1913 ( .A(n2030), .B(n2029), .C(n288), .D(n1278), .Q(n2031) );
  NAND22 U1914 ( .A(\position1/n1537 ), .B(n472), .Q(n2030) );
  AOI221 U1915 ( .A(\position1/n1340 ), .B(n603), .C(n1698), .D(n1697), .Q(
        n1699) );
  NAND22 U1916 ( .A(n261), .B(n1057), .Q(n1698) );
  AOI221 U1917 ( .A(n1696), .B(n1695), .C(n288), .D(n1059), .Q(n1697) );
  NAND22 U1918 ( .A(\position1/n1341 ), .B(n472), .Q(n1696) );
  NOR21 U1919 ( .A(n1196), .B(n43), .Q(n1922) );
  NOR21 U1920 ( .A(n604), .B(\position1/n1489 ), .Q(n1920) );
  NOR21 U1921 ( .A(n977), .B(n263), .Q(n1588) );
  NOR21 U1922 ( .A(n604), .B(\position1/n1293 ), .Q(n1586) );
  AOI221 U1923 ( .A(\position1/n1534 ), .B(n601), .C(n2036), .D(n2035), .Q(
        n2037) );
  NAND22 U1924 ( .A(n39), .B(n1272), .Q(n2036) );
  AOI221 U1925 ( .A(n2034), .B(n2033), .C(n292), .D(n1274), .Q(n2035) );
  NAND22 U1926 ( .A(\position1/n1535 ), .B(n474), .Q(n2034) );
  AOI221 U1927 ( .A(\position1/n1338 ), .B(n599), .C(n1702), .D(n1701), .Q(
        n1703) );
  NAND22 U1928 ( .A(n294), .B(n1053), .Q(n1702) );
  AOI221 U1929 ( .A(n1700), .B(n1699), .C(n292), .D(n1055), .Q(n1701) );
  NAND22 U1930 ( .A(\position1/n1339 ), .B(n474), .Q(n1700) );
  AOI221 U1931 ( .A(\position1/n1532 ), .B(n597), .C(n2040), .D(n2039), .Q(
        n2041) );
  NAND22 U1932 ( .A(n67), .B(n1268), .Q(n2040) );
  AOI221 U1933 ( .A(n2038), .B(n2037), .C(n267), .D(n1270), .Q(n2039) );
  NAND22 U1934 ( .A(\position1/n1533 ), .B(n475), .Q(n2038) );
  AOI221 U1935 ( .A(\position1/n1336 ), .B(n597), .C(n1706), .D(n1705), .Q(
        n1707) );
  NAND22 U1936 ( .A(n269), .B(n1049), .Q(n1706) );
  AOI221 U1937 ( .A(n1704), .B(n1703), .C(n296), .D(n1051), .Q(n1705) );
  NAND22 U1938 ( .A(\position1/n1337 ), .B(n475), .Q(n1704) );
  INV3 U1939 ( .A(\position1/N1659 ), .Q(n1260) );
  NOR21 U1940 ( .A(\position1/N1659 ), .B(n248), .Q(n1980) );
  INV3 U1941 ( .A(\position1/N2076 ), .Q(n1041) );
  NOR21 U1942 ( .A(\position1/N2076 ), .B(n41), .Q(n1646) );
  INV3 U1943 ( .A(\position1/N1657 ), .Q(n1262) );
  NOR21 U1944 ( .A(\position1/N1657 ), .B(n272), .Q(n1976) );
  INV3 U1945 ( .A(\position1/N2074 ), .Q(n1043) );
  NOR21 U1946 ( .A(\position1/N2074 ), .B(n245), .Q(n1642) );
  INV3 U1947 ( .A(\position1/N1661 ), .Q(n1258) );
  NOR21 U1948 ( .A(\position1/N1661 ), .B(n45), .Q(n1984) );
  INV3 U1949 ( .A(\position1/N2078 ), .Q(n1039) );
  NOR21 U1950 ( .A(\position1/N2078 ), .B(n252), .Q(n1650) );
  INV3 U1951 ( .A(\position1/N1663 ), .Q(n1256) );
  NOR21 U1952 ( .A(\position1/N1663 ), .B(n256), .Q(n1988) );
  INV3 U1953 ( .A(\position1/N2080 ), .Q(n1037) );
  NOR21 U1954 ( .A(\position1/N2080 ), .B(n40), .Q(n1654) );
  INV3 U1955 ( .A(\position1/N1665 ), .Q(n1254) );
  NOR21 U1956 ( .A(\position1/N1665 ), .B(n46), .Q(n1992) );
  INV3 U1957 ( .A(\position1/N2082 ), .Q(n1035) );
  NOR21 U1958 ( .A(\position1/N2082 ), .B(n288), .Q(n1658) );
  INV3 U1959 ( .A(\position1/N1667 ), .Q(n1252) );
  NOR21 U1960 ( .A(\position1/N1667 ), .B(n43), .Q(n1996) );
  INV3 U1961 ( .A(\position1/N2084 ), .Q(n1033) );
  NOR21 U1962 ( .A(\position1/N2084 ), .B(n292), .Q(n1662) );
  INV3 U1963 ( .A(\position1/N1669 ), .Q(n1250) );
  NOR21 U1964 ( .A(\position1/N1669 ), .B(n42), .Q(n2000) );
  INV3 U1965 ( .A(\position1/N2086 ), .Q(n1031) );
  NOR21 U1966 ( .A(\position1/N2086 ), .B(n296), .Q(n1666) );
  AOI221 U1967 ( .A(n2046), .B(n2045), .C(n516), .D(n1302), .Q(n2047) );
  INV3 U1968 ( .A(\position1/N1553 ), .Q(n1302) );
  NOR31 U1969 ( .A(\position1/N1573 ), .B(\position1/N1548 ), .C(
        \position1/N1547 ), .Q(n2046) );
  NOR40 U1970 ( .A(\position1/N1552 ), .B(\position1/N1551 ), .C(
        \position1/N1550 ), .D(\position1/N1549 ), .Q(n2045) );
  AOI221 U1971 ( .A(n1712), .B(n1711), .C(n516), .D(n1083), .Q(n1713) );
  INV3 U1972 ( .A(\position1/N1970 ), .Q(n1083) );
  NOR31 U1973 ( .A(\position1/N1990 ), .B(\position1/N1965 ), .C(
        \position1/N1964 ), .Q(n1712) );
  NOR40 U1974 ( .A(\position1/N1969 ), .B(\position1/N1968 ), .C(
        \position1/N1967 ), .D(\position1/N1966 ), .Q(n1711) );
  AOI221 U1975 ( .A(n1166), .B(n269), .C(n1888), .D(n1887), .Q(n1889) );
  NAND22 U1976 ( .A(n598), .B(\position1/n1461 ), .Q(n1887) );
  AOI221 U1977 ( .A(n1886), .B(n1885), .C(n475), .D(\position1/n1462 ), .Q(
        n1888) );
  AOI221 U1978 ( .A(n947), .B(n298), .C(n1554), .D(n1553), .Q(n1555) );
  NAND22 U1979 ( .A(n598), .B(\position1/n1265 ), .Q(n1553) );
  AOI221 U1980 ( .A(n1552), .B(n1551), .C(\position1/N2447 ), .D(
        \position1/n1266 ), .Q(n1554) );
  AOI2111 U1981 ( .A(n1144), .B(n256), .C(n1839), .D(n1145), .Q(n1840) );
  INV3 U1982 ( .A(n1838), .Q(n1145) );
  NOR21 U1983 ( .A(n614), .B(\position1/n1445 ), .Q(n1839) );
  OAI2111 U1984 ( .A(n280), .B(n1147), .C(n1837), .D(n1836), .Q(n1838) );
  AOI2111 U1985 ( .A(n925), .B(n284), .C(n1505), .D(n926), .Q(n1506) );
  INV3 U1986 ( .A(n1504), .Q(n926) );
  NOR21 U1987 ( .A(n613), .B(\position1/n1249 ), .Q(n1505) );
  OAI2111 U1988 ( .A(n252), .B(n928), .C(n1503), .D(n1502), .Q(n1504) );
  AOI221 U1989 ( .A(n1950), .B(n1949), .C(n284), .D(n1225), .Q(n1951) );
  NAND22 U1990 ( .A(\position1/n1516 ), .B(\position1/N2453 ), .Q(n1950) );
  AOI221 U1991 ( .A(\position1/n1517 ), .B(n615), .C(n1948), .D(n1947), .Q(
        n1949) );
  NAND22 U1992 ( .A(n282), .B(n1226), .Q(n1948) );
  AOI221 U1993 ( .A(n1616), .B(n1615), .C(n256), .D(n1006), .Q(n1617) );
  NAND22 U1994 ( .A(\position1/n1320 ), .B(\position1/N2453 ), .Q(n1616) );
  AOI221 U1995 ( .A(\position1/n1321 ), .B(n613), .C(n1614), .D(n1613), .Q(
        n1615) );
  NAND22 U1996 ( .A(n254), .B(n1007), .Q(n1614) );
  AOI221 U1997 ( .A(n1954), .B(n1953), .C(n259), .D(n1223), .Q(n1955) );
  NAND22 U1998 ( .A(\position1/n1514 ), .B(n472), .Q(n1954) );
  AOI221 U1999 ( .A(\position1/n1515 ), .B(n610), .C(n1952), .D(n1951), .Q(
        n1953) );
  NAND22 U2000 ( .A(n286), .B(n1224), .Q(n1952) );
  AOI221 U2001 ( .A(n1620), .B(n1619), .C(n288), .D(n1004), .Q(n1621) );
  NAND22 U2002 ( .A(\position1/n1318 ), .B(n472), .Q(n1620) );
  AOI221 U2003 ( .A(\position1/n1319 ), .B(n609), .C(n1618), .D(n1617), .Q(
        n1619) );
  NAND22 U2004 ( .A(n286), .B(n1005), .Q(n1618) );
  AOI221 U2005 ( .A(n1958), .B(n1957), .C(n263), .D(n1221), .Q(n1959) );
  NAND22 U2006 ( .A(\position1/n1512 ), .B(\position1/N2449 ), .Q(n1958) );
  AOI221 U2007 ( .A(\position1/n1513 ), .B(n605), .C(n1956), .D(n1955), .Q(
        n1957) );
  NAND22 U2008 ( .A(n38), .B(n1222), .Q(n1956) );
  AOI221 U2009 ( .A(n1624), .B(n1623), .C(n292), .D(n1002), .Q(n1625) );
  NAND22 U2010 ( .A(\position1/n1316 ), .B(\position1/N2449 ), .Q(n1624) );
  AOI221 U2011 ( .A(\position1/n1317 ), .B(n605), .C(n1622), .D(n1621), .Q(
        n1623) );
  NAND22 U2012 ( .A(n290), .B(n1003), .Q(n1622) );
  AOI221 U2013 ( .A(n1962), .B(n1961), .C(n267), .D(n1219), .Q(n1963) );
  NAND22 U2014 ( .A(\position1/n1510 ), .B(\position1/N2447 ), .Q(n1962) );
  AOI221 U2015 ( .A(\position1/n1511 ), .B(n601), .C(n1960), .D(n1959), .Q(
        n1961) );
  NAND22 U2016 ( .A(n39), .B(n1220), .Q(n1960) );
  AOI221 U2017 ( .A(n1628), .B(n1627), .C(n296), .D(n1000), .Q(n1629) );
  NAND22 U2018 ( .A(\position1/n1314 ), .B(\position1/N2447 ), .Q(n1628) );
  AOI221 U2019 ( .A(\position1/n1315 ), .B(n601), .C(n1626), .D(n1625), .Q(
        n1627) );
  NAND22 U2020 ( .A(n265), .B(n1001), .Q(n1626) );
  AOI221 U2021 ( .A(n1946), .B(n1227), .C(n280), .D(n1228), .Q(n1947) );
  INV3 U2022 ( .A(n1945), .Q(n1227) );
  NAND22 U2023 ( .A(\position1/n1519 ), .B(n619), .Q(n1946) );
  AOI221 U2024 ( .A(n1612), .B(n1008), .C(n252), .D(n1009), .Q(n1613) );
  INV3 U2025 ( .A(n1611), .Q(n1008) );
  NAND22 U2026 ( .A(\position1/n1323 ), .B(n619), .Q(n1612) );
  AOI211 U2027 ( .A(n1299), .B(n513), .C(n2011), .Q(n2012) );
  AOI221 U2028 ( .A(n2010), .B(n2009), .C(n516), .D(\position1/n1547 ), .Q(
        n2011) );
  AOI211 U2029 ( .A(n1080), .B(n34), .C(n1677), .Q(n1678) );
  AOI221 U2030 ( .A(n1676), .B(n1675), .C(n516), .D(\position1/n1351 ), .Q(
        n1677) );
  AOI221 U2031 ( .A(n2053), .B(n2052), .C(n623), .D(n1305), .Q(n2055) );
  INV3 U2032 ( .A(\position1/N1556 ), .Q(n1305) );
  NAND22 U2033 ( .A(\position1/N1556 ), .B(n246), .Q(n2052) );
  AOI221 U2034 ( .A(\position1/N1555 ), .B(n66), .C(n2051), .D(n2050), .Q(
        n2053) );
  AOI221 U2035 ( .A(n1719), .B(n1718), .C(n623), .D(n1086), .Q(n1721) );
  INV3 U2036 ( .A(\position1/N1973 ), .Q(n1086) );
  NAND22 U2037 ( .A(\position1/N1973 ), .B(n246), .Q(n1718) );
  AOI221 U2038 ( .A(\position1/N1972 ), .B(n245), .C(n1717), .D(n1716), .Q(
        n1719) );
  AOI221 U2039 ( .A(n1174), .B(n282), .C(n1872), .D(n1871), .Q(n1874) );
  NAND22 U2040 ( .A(n615), .B(\position1/n1469 ), .Q(n1871) );
  AOI221 U2041 ( .A(n1870), .B(n1869), .C(n469), .D(\position1/n1470 ), .Q(
        n1872) );
  NAND22 U2042 ( .A(n1175), .B(n45), .Q(n1869) );
  AOI221 U2043 ( .A(n955), .B(n254), .C(n1538), .D(n1537), .Q(n1540) );
  NAND22 U2044 ( .A(n615), .B(\position1/n1273 ), .Q(n1537) );
  AOI221 U2045 ( .A(n1536), .B(n1535), .C(n470), .D(\position1/n1274 ), .Q(
        n1538) );
  NAND22 U2046 ( .A(n956), .B(n45), .Q(n1535) );
  AOI221 U2047 ( .A(n2057), .B(n2056), .C(n620), .D(n1307), .Q(n2059) );
  INV3 U2048 ( .A(\position1/N1558 ), .Q(n1307) );
  NAND22 U2049 ( .A(\position1/N1558 ), .B(n250), .Q(n2056) );
  AOI221 U2050 ( .A(\position1/N1557 ), .B(n248), .C(n2055), .D(n2054), .Q(
        n2057) );
  AOI221 U2051 ( .A(n1723), .B(n1722), .C(n620), .D(n1088), .Q(n1725) );
  INV3 U2052 ( .A(\position1/N1975 ), .Q(n1088) );
  NAND22 U2053 ( .A(\position1/N1975 ), .B(n250), .Q(n1722) );
  AOI221 U2054 ( .A(\position1/N1974 ), .B(n41), .C(n1721), .D(n1720), .Q(
        n1723) );
  AOI221 U2055 ( .A(n2061), .B(n2060), .C(n616), .D(n1309), .Q(n2063) );
  INV3 U2056 ( .A(\position1/N1560 ), .Q(n1309) );
  NAND22 U2057 ( .A(\position1/N1560 ), .B(n100), .Q(n2060) );
  AOI221 U2058 ( .A(\position1/N1559 ), .B(n252), .C(n2059), .D(n2058), .Q(
        n2061) );
  AOI221 U2059 ( .A(n1727), .B(n1726), .C(n612), .D(n1090), .Q(n1729) );
  INV3 U2060 ( .A(\position1/N1977 ), .Q(n1090) );
  NAND22 U2061 ( .A(\position1/N1977 ), .B(n282), .Q(n1726) );
  AOI221 U2062 ( .A(\position1/N1976 ), .B(n252), .C(n1725), .D(n1724), .Q(
        n1727) );
  AOI221 U2063 ( .A(n2065), .B(n2064), .C(n611), .D(n1311), .Q(n2067) );
  INV3 U2064 ( .A(\position1/N1562 ), .Q(n1311) );
  NAND22 U2065 ( .A(\position1/N1562 ), .B(n286), .Q(n2064) );
  AOI221 U2066 ( .A(\position1/N1561 ), .B(n256), .C(n2063), .D(n2062), .Q(
        n2065) );
  AOI221 U2067 ( .A(n1731), .B(n1730), .C(n610), .D(n1092), .Q(n1733) );
  INV3 U2068 ( .A(\position1/N1979 ), .Q(n1092) );
  NAND22 U2069 ( .A(\position1/N1979 ), .B(n286), .Q(n1730) );
  AOI221 U2070 ( .A(\position1/N1978 ), .B(n284), .C(n1729), .D(n1728), .Q(
        n1731) );
  AOI221 U2071 ( .A(n2069), .B(n2068), .C(n606), .D(n1313), .Q(n2071) );
  INV3 U2072 ( .A(\position1/N1564 ), .Q(n1313) );
  NAND22 U2073 ( .A(\position1/N1564 ), .B(n38), .Q(n2068) );
  AOI221 U2074 ( .A(\position1/N1563 ), .B(n259), .C(n2067), .D(n2066), .Q(
        n2069) );
  AOI221 U2075 ( .A(n1735), .B(n1734), .C(n606), .D(n1094), .Q(n1737) );
  INV3 U2076 ( .A(\position1/N1981 ), .Q(n1094) );
  NAND22 U2077 ( .A(\position1/N1981 ), .B(n290), .Q(n1734) );
  AOI221 U2078 ( .A(\position1/N1980 ), .B(n259), .C(n1733), .D(n1732), .Q(
        n1735) );
  AOI221 U2079 ( .A(n2073), .B(n2072), .C(n602), .D(n1315), .Q(n2075) );
  INV3 U2080 ( .A(\position1/N1566 ), .Q(n1315) );
  NAND22 U2081 ( .A(\position1/N1566 ), .B(n39), .Q(n2072) );
  AOI221 U2082 ( .A(\position1/N1565 ), .B(n263), .C(n2071), .D(n2070), .Q(
        n2073) );
  AOI221 U2083 ( .A(n1739), .B(n1738), .C(n602), .D(n1096), .Q(n1741) );
  INV3 U2084 ( .A(\position1/N1983 ), .Q(n1096) );
  NAND22 U2085 ( .A(\position1/N1983 ), .B(n294), .Q(n1738) );
  AOI221 U2086 ( .A(\position1/N1982 ), .B(n43), .C(n1737), .D(n1736), .Q(
        n1739) );
  AOI221 U2087 ( .A(n2077), .B(n2076), .C(n598), .D(n1317), .Q(n2079) );
  INV3 U2088 ( .A(\position1/N1568 ), .Q(n1317) );
  NAND22 U2089 ( .A(\position1/N1568 ), .B(n67), .Q(n2076) );
  AOI221 U2090 ( .A(\position1/N1567 ), .B(n267), .C(n2075), .D(n2074), .Q(
        n2077) );
  AOI221 U2091 ( .A(n1743), .B(n1742), .C(n598), .D(n1098), .Q(n1745) );
  INV3 U2092 ( .A(\position1/N1985 ), .Q(n1098) );
  NAND22 U2093 ( .A(\position1/N1985 ), .B(n298), .Q(n1742) );
  AOI221 U2094 ( .A(\position1/N1984 ), .B(n42), .C(n1741), .D(n1740), .Q(
        n1743) );
  AOI221 U2095 ( .A(n1804), .B(n1803), .C(n606), .D(\position1/n1417 ), .Q(
        n1806) );
  NAND22 U2096 ( .A(n1110), .B(n261), .Q(n1803) );
  AOI221 U2097 ( .A(n1112), .B(n288), .C(n1111), .D(n1802), .Q(n1804) );
  INV3 U2098 ( .A(\position1/n1417 ), .Q(n1110) );
  AOI221 U2099 ( .A(n1470), .B(n1469), .C(n606), .D(\position1/n1221 ), .Q(
        n1472) );
  NAND22 U2100 ( .A(n891), .B(n290), .Q(n1469) );
  AOI221 U2101 ( .A(n893), .B(n259), .C(n892), .D(n1468), .Q(n1470) );
  INV3 U2102 ( .A(\position1/n1221 ), .Q(n891) );
  AOI221 U2103 ( .A(n1808), .B(n1807), .C(n602), .D(\position1/n1415 ), .Q(
        n1810) );
  NAND22 U2104 ( .A(n1108), .B(n294), .Q(n1807) );
  AOI221 U2105 ( .A(n1109), .B(n43), .C(n1806), .D(n1805), .Q(n1808) );
  INV3 U2106 ( .A(\position1/n1415 ), .Q(n1108) );
  AOI221 U2107 ( .A(n1474), .B(n1473), .C(n602), .D(\position1/n1219 ), .Q(
        n1476) );
  NAND22 U2108 ( .A(n889), .B(n265), .Q(n1473) );
  AOI221 U2109 ( .A(n890), .B(n263), .C(n1472), .D(n1471), .Q(n1474) );
  INV3 U2110 ( .A(\position1/n1219 ), .Q(n889) );
  AOI221 U2111 ( .A(n1812), .B(n1811), .C(n598), .D(\position1/n1413 ), .Q(
        n1814) );
  NAND22 U2112 ( .A(n1106), .B(n269), .Q(n1811) );
  AOI221 U2113 ( .A(n1107), .B(n42), .C(n1810), .D(n1809), .Q(n1812) );
  INV3 U2114 ( .A(\position1/n1413 ), .Q(n1106) );
  AOI221 U2115 ( .A(n1478), .B(n1477), .C(n598), .D(\position1/n1217 ), .Q(
        n1480) );
  NAND22 U2116 ( .A(n887), .B(n298), .Q(n1477) );
  AOI221 U2117 ( .A(n888), .B(n267), .C(n1476), .D(n1475), .Q(n1478) );
  INV3 U2118 ( .A(\position1/n1217 ), .Q(n887) );
  AOI221 U2119 ( .A(n1178), .B(n274), .C(n1864), .D(n1863), .Q(n1866) );
  NAND22 U2120 ( .A(n622), .B(\position1/n1473 ), .Q(n1863) );
  AOI221 U2121 ( .A(n1862), .B(n1861), .C(n627), .D(\position1/n1474 ), .Q(
        n1864) );
  NAND22 U2122 ( .A(n1179), .B(n66), .Q(n1861) );
  AOI221 U2123 ( .A(n959), .B(n274), .C(n1530), .D(n1529), .Q(n1532) );
  NAND22 U2124 ( .A(n623), .B(\position1/n1277 ), .Q(n1529) );
  AOI221 U2125 ( .A(n1528), .B(n1527), .C(n627), .D(\position1/n1278 ), .Q(
        n1530) );
  NAND22 U2126 ( .A(n960), .B(n272), .Q(n1527) );
  AOI221 U2127 ( .A(n1176), .B(n278), .C(n1868), .D(n1867), .Q(n1870) );
  NAND22 U2128 ( .A(n620), .B(\position1/n1471 ), .Q(n1867) );
  AOI221 U2129 ( .A(n1866), .B(n1865), .C(n468), .D(\position1/n1472 ), .Q(
        n1868) );
  NAND22 U2130 ( .A(n1177), .B(n41), .Q(n1865) );
  AOI221 U2131 ( .A(n957), .B(n250), .C(n1534), .D(n1533), .Q(n1536) );
  NAND22 U2132 ( .A(n620), .B(\position1/n1275 ), .Q(n1533) );
  AOI221 U2133 ( .A(n1532), .B(n1531), .C(\position1/N2457 ), .D(
        \position1/n1276 ), .Q(n1534) );
  NAND22 U2134 ( .A(n958), .B(n248), .Q(n1531) );
  AOI221 U2135 ( .A(n1170), .B(n261), .C(n1880), .D(n1879), .Q(n1882) );
  NAND22 U2136 ( .A(n605), .B(\position1/n1465 ), .Q(n1879) );
  AOI221 U2137 ( .A(n1878), .B(n1877), .C(n473), .D(\position1/n1466 ), .Q(
        n1880) );
  NAND22 U2138 ( .A(n1171), .B(n46), .Q(n1877) );
  AOI221 U2139 ( .A(n951), .B(n290), .C(n1546), .D(n1545), .Q(n1548) );
  NAND22 U2140 ( .A(n605), .B(\position1/n1269 ), .Q(n1545) );
  AOI221 U2141 ( .A(n1544), .B(n1543), .C(n473), .D(\position1/n1270 ), .Q(
        n1546) );
  NAND22 U2142 ( .A(n952), .B(n46), .Q(n1543) );
  AOI221 U2143 ( .A(n1168), .B(n294), .C(n1884), .D(n1883), .Q(n1886) );
  NAND22 U2144 ( .A(n601), .B(\position1/n1463 ), .Q(n1883) );
  AOI221 U2145 ( .A(n1882), .B(n1881), .C(n474), .D(\position1/n1464 ), .Q(
        n1884) );
  NAND22 U2146 ( .A(n1169), .B(n43), .Q(n1881) );
  AOI221 U2147 ( .A(n949), .B(n265), .C(n1550), .D(n1549), .Q(n1552) );
  NAND22 U2148 ( .A(n601), .B(\position1/n1267 ), .Q(n1549) );
  AOI221 U2149 ( .A(n1548), .B(n1547), .C(\position1/N2449 ), .D(
        \position1/n1268 ), .Q(n1550) );
  NAND22 U2150 ( .A(n950), .B(n43), .Q(n1547) );
  AOI221 U2151 ( .A(n1180), .B(n273), .C(n1860), .D(n1859), .Q(n1862) );
  NAND22 U2152 ( .A(n631), .B(\position1/n1475 ), .Q(n1859) );
  AOI211 U2153 ( .A(n517), .B(\position1/n1476 ), .C(n1858), .Q(n1860) );
  AOI2111 U2154 ( .A(n1181), .B(n34), .C(n1182), .D(n1183), .Q(n1858) );
  AOI221 U2155 ( .A(n961), .B(n273), .C(n1526), .D(n1525), .Q(n1528) );
  NAND22 U2156 ( .A(n631), .B(\position1/n1279 ), .Q(n1525) );
  AOI211 U2157 ( .A(n517), .B(\position1/n1280 ), .C(n1524), .Q(n1526) );
  AOI2111 U2158 ( .A(n962), .B(n34), .C(n963), .D(n964), .Q(n1524) );
  AOI221 U2159 ( .A(n1172), .B(n286), .C(n1876), .D(n1875), .Q(n1878) );
  NAND22 U2160 ( .A(n610), .B(\position1/n1467 ), .Q(n1875) );
  AOI221 U2161 ( .A(n1874), .B(n1873), .C(n471), .D(\position1/n1468 ), .Q(
        n1876) );
  NAND22 U2162 ( .A(n1173), .B(n40), .Q(n1873) );
  AOI221 U2163 ( .A(n953), .B(n286), .C(n1542), .D(n1541), .Q(n1544) );
  NAND22 U2164 ( .A(n610), .B(\position1/n1271 ), .Q(n1541) );
  AOI221 U2165 ( .A(n1540), .B(n1539), .C(\position1/N2453 ), .D(
        \position1/n1272 ), .Q(n1542) );
  NAND22 U2166 ( .A(n954), .B(n256), .Q(n1539) );
  AOI221 U2167 ( .A(n1788), .B(n1787), .C(n623), .D(\position1/n1425 ), .Q(
        n1790) );
  NAND22 U2168 ( .A(n1119), .B(n274), .Q(n1787) );
  AOI221 U2169 ( .A(n1120), .B(n272), .C(n1786), .D(n1785), .Q(n1788) );
  INV3 U2170 ( .A(\position1/n1425 ), .Q(n1119) );
  AOI221 U2171 ( .A(n1454), .B(n1453), .C(n623), .D(\position1/n1229 ), .Q(
        n1456) );
  NAND22 U2172 ( .A(n900), .B(n246), .Q(n1453) );
  AOI221 U2173 ( .A(n901), .B(n245), .C(n1452), .D(n1451), .Q(n1454) );
  INV3 U2174 ( .A(\position1/n1229 ), .Q(n900) );
  AOI221 U2175 ( .A(n1792), .B(n1791), .C(n620), .D(\position1/n1423 ), .Q(
        n1794) );
  NAND22 U2176 ( .A(n1117), .B(n278), .Q(n1791) );
  AOI221 U2177 ( .A(n1118), .B(n276), .C(n1790), .D(n1789), .Q(n1792) );
  INV3 U2178 ( .A(\position1/n1423 ), .Q(n1117) );
  AOI221 U2179 ( .A(n1458), .B(n1457), .C(n620), .D(\position1/n1227 ), .Q(
        n1460) );
  NAND22 U2180 ( .A(n898), .B(n250), .Q(n1457) );
  AOI221 U2181 ( .A(n899), .B(n248), .C(n1456), .D(n1455), .Q(n1458) );
  INV3 U2182 ( .A(\position1/n1227 ), .Q(n898) );
  AOI221 U2183 ( .A(n2049), .B(n2048), .C(n632), .D(n1303), .Q(n2051) );
  INV3 U2184 ( .A(\position1/N1554 ), .Q(n1303) );
  NAND22 U2185 ( .A(\position1/N1554 ), .B(n628), .Q(n2048) );
  AOI211 U2186 ( .A(\position1/N1553 ), .B(n513), .C(n2047), .Q(n2049) );
  AOI221 U2187 ( .A(n1715), .B(n1714), .C(n632), .D(n1084), .Q(n1717) );
  INV3 U2188 ( .A(\position1/N1971 ), .Q(n1084) );
  NAND22 U2189 ( .A(\position1/N1971 ), .B(n273), .Q(n1714) );
  AOI211 U2190 ( .A(\position1/N1970 ), .B(n34), .C(n1713), .Q(n1715) );
  INV3 U2191 ( .A(\position1/N1656 ), .Q(n1263) );
  AOI211 U2192 ( .A(\position1/N1655 ), .B(n513), .C(n1972), .Q(n1973) );
  AOI221 U2193 ( .A(n1971), .B(n1970), .C(n516), .D(n1264), .Q(n1972) );
  INV3 U2194 ( .A(\position1/N2073 ), .Q(n1044) );
  AOI211 U2195 ( .A(\position1/N2072 ), .B(n34), .C(n1638), .Q(n1639) );
  AOI221 U2196 ( .A(n1637), .B(n1636), .C(n516), .D(n1045), .Q(n1638) );
  INV3 U2197 ( .A(n166), .Q(\position1/sub_216_I2/carry [8]) );
  NOR21 U2198 ( .A(n513), .B(\position1/N1553 ), .Q(n166) );
  INV3 U2199 ( .A(n172), .Q(\position1/sub_226_I2/carry [8]) );
  NOR21 U2200 ( .A(n513), .B(\position1/N1970 ), .Q(n172) );
  INV3 U2201 ( .A(\position1/N1519 ), .Q(n521) );
  INV3 U2202 ( .A(\position1/N1936 ), .Q(n555) );
  AOI211 U2203 ( .A(n632), .B(n1784), .C(n1121), .Q(n1786) );
  INV3 U2204 ( .A(n1783), .Q(n1121) );
  NAND22 U2205 ( .A(n1122), .B(n34), .Q(n1784) );
  AOI211 U2206 ( .A(n632), .B(n1450), .C(n902), .Q(n1452) );
  INV3 U2207 ( .A(n1449), .Q(n902) );
  NAND22 U2208 ( .A(n903), .B(n34), .Q(n1450) );
  NAND22 U2209 ( .A(\position1/n1545 ), .B(n625), .Q(n2008) );
  NAND22 U2210 ( .A(\position1/n1349 ), .B(n625), .Q(n1674) );
  NAND22 U2211 ( .A(\position1/n1544 ), .B(n622), .Q(n2018) );
  NAND22 U2212 ( .A(\position1/n1348 ), .B(n622), .Q(n1684) );
  NOR21 U2213 ( .A(n618), .B(\position1/n1519 ), .Q(n1944) );
  NOR21 U2214 ( .A(n619), .B(\position1/n1323 ), .Q(n1610) );
  BUF2 U2215 ( .A(\position1/n1152 ), .Q(n485) );
  NAND22 U2216 ( .A(n594), .B(\position1/n1460 ), .Q(n1892) );
  NAND22 U2217 ( .A(n593), .B(\position1/n1264 ), .Q(n1558) );
  NOR21 U2218 ( .A(n51), .B(n630), .Q(n2084) );
  NOR21 U2219 ( .A(n50), .B(n630), .Q(n1750) );
  BUF2 U2220 ( .A(n101), .Q(n589) );
  BUF2 U2221 ( .A(n590), .Q(n588) );
  NAND22 U2222 ( .A(n610), .B(\position1/n1419 ), .Q(n1802) );
  NAND22 U2223 ( .A(n610), .B(\position1/n1223 ), .Q(n1468) );
  NAND22 U2224 ( .A(\position1/N2449 ), .B(\position1/n1416 ), .Q(n1805) );
  NAND22 U2225 ( .A(\position1/N2449 ), .B(\position1/n1220 ), .Q(n1471) );
  NAND22 U2226 ( .A(\position1/N2447 ), .B(\position1/n1414 ), .Q(n1809) );
  NAND22 U2227 ( .A(\position1/N2447 ), .B(\position1/n1218 ), .Q(n1475) );
  NAND22 U2228 ( .A(n593), .B(\position1/n1412 ), .Q(n1813) );
  NAND22 U2229 ( .A(n594), .B(\position1/n1216 ), .Q(n1479) );
  NAND22 U2230 ( .A(n627), .B(\position1/n1426 ), .Q(n1785) );
  NAND22 U2231 ( .A(n627), .B(\position1/n1230 ), .Q(n1451) );
  NAND22 U2232 ( .A(\position1/N2457 ), .B(\position1/n1424 ), .Q(n1789) );
  NAND22 U2233 ( .A(\position1/N2457 ), .B(\position1/n1228 ), .Q(n1455) );
  NAND22 U2234 ( .A(n470), .B(\position1/n1422 ), .Q(n1793) );
  NAND22 U2235 ( .A(n470), .B(\position1/n1226 ), .Q(n1459) );
  NAND22 U2236 ( .A(\position1/n1445 ), .B(n614), .Q(n1837) );
  NAND22 U2237 ( .A(\position1/n1249 ), .B(n614), .Q(n1503) );
  NAND22 U2238 ( .A(\position1/n1531 ), .B(n592), .Q(n2042) );
  NAND22 U2239 ( .A(\position1/n1335 ), .B(n592), .Q(n1708) );
  NOR21 U2240 ( .A(n600), .B(\position1/n1487 ), .Q(n1924) );
  NOR21 U2241 ( .A(n600), .B(\position1/n1291 ), .Q(n1590) );
  NOR21 U2242 ( .A(n622), .B(n1261), .Q(n1978) );
  INV3 U2243 ( .A(\position1/N1658 ), .Q(n1261) );
  NOR21 U2244 ( .A(n621), .B(n1042), .Q(n1644) );
  INV3 U2245 ( .A(\position1/N2075 ), .Q(n1042) );
  NOR21 U2246 ( .A(n613), .B(n1257), .Q(n1986) );
  INV3 U2247 ( .A(\position1/N1662 ), .Q(n1257) );
  NOR21 U2248 ( .A(n614), .B(n1038), .Q(n1652) );
  INV3 U2249 ( .A(\position1/N2079 ), .Q(n1038) );
  NOR21 U2250 ( .A(n608), .B(n1255), .Q(n1990) );
  INV3 U2251 ( .A(\position1/N1664 ), .Q(n1255) );
  NOR21 U2252 ( .A(n608), .B(n1036), .Q(n1656) );
  INV3 U2253 ( .A(\position1/N2081 ), .Q(n1036) );
  NOR21 U2254 ( .A(n604), .B(n1253), .Q(n1994) );
  INV3 U2255 ( .A(\position1/N1666 ), .Q(n1253) );
  NOR21 U2256 ( .A(n604), .B(n1034), .Q(n1660) );
  INV3 U2257 ( .A(\position1/N2083 ), .Q(n1034) );
  NOR21 U2258 ( .A(n600), .B(n1251), .Q(n1998) );
  INV3 U2259 ( .A(\position1/N1668 ), .Q(n1251) );
  NOR21 U2260 ( .A(n600), .B(n1032), .Q(n1664) );
  INV3 U2261 ( .A(\position1/N2085 ), .Q(n1032) );
  NOR21 U2262 ( .A(n596), .B(n1249), .Q(n2002) );
  INV3 U2263 ( .A(\position1/N1670 ), .Q(n1249) );
  NOR21 U2264 ( .A(n596), .B(n1030), .Q(n1668) );
  INV3 U2265 ( .A(\position1/N2087 ), .Q(n1030) );
  NOR21 U2266 ( .A(n618), .B(n1259), .Q(n1982) );
  INV3 U2267 ( .A(\position1/N1660 ), .Q(n1259) );
  NOR21 U2268 ( .A(n618), .B(n1040), .Q(n1648) );
  INV3 U2269 ( .A(\position1/N2077 ), .Q(n1040) );
  NAND22 U2270 ( .A(n627), .B(n1304), .Q(n2050) );
  INV3 U2271 ( .A(\position1/N1555 ), .Q(n1304) );
  NAND22 U2272 ( .A(n626), .B(n1085), .Q(n1716) );
  INV3 U2273 ( .A(\position1/N1972 ), .Q(n1085) );
  NAND22 U2274 ( .A(n468), .B(n1306), .Q(n2054) );
  INV3 U2275 ( .A(\position1/N1557 ), .Q(n1306) );
  NAND22 U2276 ( .A(n468), .B(n1087), .Q(n1720) );
  INV3 U2277 ( .A(\position1/N1974 ), .Q(n1087) );
  NAND22 U2278 ( .A(n469), .B(n1308), .Q(n2058) );
  INV3 U2279 ( .A(\position1/N1559 ), .Q(n1308) );
  NAND22 U2280 ( .A(n469), .B(n1089), .Q(n1724) );
  INV3 U2281 ( .A(\position1/N1976 ), .Q(n1089) );
  NAND22 U2282 ( .A(n471), .B(n1310), .Q(n2062) );
  INV3 U2283 ( .A(\position1/N1561 ), .Q(n1310) );
  NAND22 U2284 ( .A(n471), .B(n1091), .Q(n1728) );
  INV3 U2285 ( .A(\position1/N1978 ), .Q(n1091) );
  NAND22 U2286 ( .A(n473), .B(n1312), .Q(n2066) );
  INV3 U2287 ( .A(\position1/N1563 ), .Q(n1312) );
  NAND22 U2288 ( .A(n473), .B(n1093), .Q(n1732) );
  INV3 U2289 ( .A(\position1/N1980 ), .Q(n1093) );
  NAND22 U2290 ( .A(n474), .B(n1314), .Q(n2070) );
  INV3 U2291 ( .A(\position1/N1565 ), .Q(n1314) );
  NAND22 U2292 ( .A(n474), .B(n1095), .Q(n1736) );
  INV3 U2293 ( .A(\position1/N1982 ), .Q(n1095) );
  NAND22 U2294 ( .A(n475), .B(n1316), .Q(n2074) );
  INV3 U2295 ( .A(\position1/N1567 ), .Q(n1316) );
  NAND22 U2296 ( .A(n475), .B(n1097), .Q(n1740) );
  INV3 U2297 ( .A(\position1/N1984 ), .Q(n1097) );
  INV3 U2298 ( .A(n1844), .Q(n1141) );
  AOI2111 U2299 ( .A(n1142), .B(n46), .C(n1843), .D(n1842), .Q(n1844) );
  NOR21 U2300 ( .A(n608), .B(\position1/n1443 ), .Q(n1843) );
  AOI2111 U2301 ( .A(n609), .B(\position1/n1443 ), .C(n1841), .D(n1840), .Q(
        n1842) );
  INV3 U2302 ( .A(n1510), .Q(n922) );
  AOI2111 U2303 ( .A(n923), .B(n259), .C(n1509), .D(n1508), .Q(n1510) );
  NOR21 U2304 ( .A(n608), .B(\position1/n1247 ), .Q(n1509) );
  AOI2111 U2305 ( .A(n609), .B(\position1/n1247 ), .C(n1507), .D(n1506), .Q(
        n1508) );
  INV3 U2306 ( .A(n1927), .Q(n1193) );
  NOR21 U2307 ( .A(n1194), .B(n42), .Q(n1926) );
  INV3 U2308 ( .A(n1593), .Q(n974) );
  NOR21 U2309 ( .A(n975), .B(n267), .Q(n1592) );
  INV3 U2310 ( .A(n1797), .Q(n1114) );
  AOI221 U2311 ( .A(n1796), .B(n1795), .C(n616), .D(\position1/n1421 ), .Q(
        n1797) );
  NAND22 U2312 ( .A(n1115), .B(n254), .Q(n1795) );
  AOI221 U2313 ( .A(n1116), .B(n45), .C(n1794), .D(n1793), .Q(n1796) );
  INV3 U2314 ( .A(n1463), .Q(n895) );
  AOI221 U2315 ( .A(n1462), .B(n1461), .C(n616), .D(\position1/n1225 ), .Q(
        n1463) );
  NAND22 U2316 ( .A(n896), .B(n282), .Q(n1461) );
  AOI221 U2317 ( .A(n897), .B(n252), .C(n1460), .D(n1459), .Q(n1462) );
  INV3 U2318 ( .A(n1801), .Q(n1111) );
  NOR21 U2319 ( .A(\position1/n1419 ), .B(n609), .Q(n1799) );
  INV3 U2320 ( .A(n1467), .Q(n892) );
  NOR21 U2321 ( .A(\position1/n1223 ), .B(n609), .Q(n1465) );
  INV3 U2322 ( .A(n2088), .Q(n1342) );
  NOR21 U2323 ( .A(n65), .B(n622), .Q(n2088) );
  INV3 U2324 ( .A(n1754), .Q(n1341) );
  NOR21 U2325 ( .A(n58), .B(n622), .Q(n1754) );
  INV3 U2326 ( .A(n2092), .Q(n1338) );
  NOR21 U2327 ( .A(n64), .B(n619), .Q(n2092) );
  INV3 U2328 ( .A(n1758), .Q(n1337) );
  NOR21 U2329 ( .A(n57), .B(n619), .Q(n1758) );
  INV3 U2330 ( .A(n2096), .Q(n1334) );
  NOR21 U2331 ( .A(n63), .B(n614), .Q(n2096) );
  INV3 U2332 ( .A(n1762), .Q(n1333) );
  NOR21 U2333 ( .A(n56), .B(n615), .Q(n1762) );
  INV3 U2334 ( .A(n2100), .Q(n1330) );
  NOR21 U2335 ( .A(n62), .B(n609), .Q(n2100) );
  INV3 U2336 ( .A(n1766), .Q(n1329) );
  NOR21 U2337 ( .A(n55), .B(n609), .Q(n1766) );
  INV3 U2338 ( .A(n2104), .Q(n1326) );
  NOR21 U2339 ( .A(n61), .B(n605), .Q(n2104) );
  INV3 U2340 ( .A(n1770), .Q(n1325) );
  NOR21 U2341 ( .A(n54), .B(n605), .Q(n1770) );
  INV3 U2342 ( .A(n2108), .Q(n1322) );
  NOR21 U2343 ( .A(n60), .B(n601), .Q(n2108) );
  INV3 U2344 ( .A(n1774), .Q(n1321) );
  NOR21 U2345 ( .A(n53), .B(n601), .Q(n1774) );
  INV3 U2346 ( .A(n2112), .Q(n1318) );
  NOR21 U2347 ( .A(n59), .B(n597), .Q(n2112) );
  INV3 U2348 ( .A(n1778), .Q(n1099) );
  NOR21 U2349 ( .A(n52), .B(n597), .Q(n1778) );
  INV3 U2350 ( .A(n1896), .Q(n1184) );
  NOR21 U2351 ( .A(n596), .B(\position1/n1485 ), .Q(n1896) );
  INV3 U2352 ( .A(n1562), .Q(n965) );
  NOR21 U2353 ( .A(n596), .B(\position1/n1289 ), .Q(n1562) );
  INV3 U2354 ( .A(n1798), .Q(n1113) );
  NAND22 U2355 ( .A(\position1/N2453 ), .B(\position1/n1420 ), .Q(n1798) );
  INV3 U2356 ( .A(n1464), .Q(n894) );
  NAND22 U2357 ( .A(\position1/N2453 ), .B(\position1/n1224 ), .Q(n1464) );
  BUF2 U2358 ( .A(n101), .Q(n590) );
  NOR40 U2359 ( .A(n816), .B(n825), .C(\gensync1/N167 ), .D(\gensync1/N168 ), 
        .Q(\gensync1/N129 ) );
  INV3 U2360 ( .A(n1371), .Q(n825) );
  INV3 U2361 ( .A(n1370), .Q(n816) );
  NOR31 U2362 ( .A(\gensync1/N166 ), .B(\gensync1/comptY[9] ), .C(
        \gensync1/N165 ), .Q(n1371) );
  NOR40 U2363 ( .A(\gensync1/N169 ), .B(\gensync1/N170 ), .C(\gensync1/N171 ), 
        .D(\gensync1/N172 ), .Q(n1370) );
  AOI211 U2364 ( .A(\gensync1/N175 ), .B(n1379), .C(\gensync1/N174 ), .Q(
        \gensync1/N72 ) );
  NAND31 U2365 ( .A(n1378), .B(n7), .C(n1377), .Q(n1379) );
  NOR31 U2366 ( .A(\gensync1/N178 ), .B(\gensync1/N176 ), .C(\gensync1/N177 ), 
        .Q(n1377) );
  NAND22 U2367 ( .A(n814), .B(n3), .Q(\gensync1/n99 ) );
  NAND41 U2368 ( .A(\position1/n860 ), .B(\position1/n861 ), .C(
        \position1/n862 ), .D(\position1/n863 ), .Q(\position1/n1587 ) );
  NAND22 U2369 ( .A(\position1/y_sum [23]), .B(n510), .Q(\position1/n861 ) );
  NAND22 U2370 ( .A(\position1/N1225 ), .B(n638), .Q(\position1/n863 ) );
  AOI221 U2371 ( .A(\position1/N558 ), .B(n512), .C(\position1/N1002 ), .D(
        n641), .Q(\position1/n862 ) );
  NAND41 U2372 ( .A(\position1/n960 ), .B(\position1/n961 ), .C(
        \position1/n962 ), .D(\position1/n963 ), .Q(\position1/n1612 ) );
  NAND22 U2373 ( .A(\position1/x_sum [23]), .B(n508), .Q(\position1/n961 ) );
  NAND22 U2374 ( .A(\position1/N1200 ), .B(n635), .Q(\position1/n963 ) );
  AOI221 U2375 ( .A(\position1/N508 ), .B(n511), .C(\position1/N927 ), .D(n639), .Q(\position1/n962 ) );
  NAND41 U2376 ( .A(\position1/n964 ), .B(\position1/n965 ), .C(
        \position1/n966 ), .D(\position1/n967 ), .Q(\position1/n1613 ) );
  NAND22 U2377 ( .A(\position1/x_sum [22]), .B(n508), .Q(\position1/n965 ) );
  NAND22 U2378 ( .A(\position1/N1199 ), .B(n635), .Q(\position1/n967 ) );
  AOI221 U2379 ( .A(\position1/N507 ), .B(n511), .C(\position1/N926 ), .D(n639), .Q(\position1/n966 ) );
  NAND41 U2380 ( .A(\position1/n852 ), .B(\position1/n853 ), .C(
        \position1/n854 ), .D(\position1/n855 ), .Q(\position1/n1586 ) );
  NAND22 U2381 ( .A(\position1/y_sum [24]), .B(n510), .Q(\position1/n853 ) );
  NAND22 U2382 ( .A(\position1/N1226 ), .B(n638), .Q(\position1/n855 ) );
  AOI221 U2383 ( .A(\position1/N559 ), .B(n512), .C(\position1/N1003 ), .D(
        n641), .Q(\position1/n854 ) );
  NAND41 U2384 ( .A(\position1/n956 ), .B(\position1/n957 ), .C(
        \position1/n958 ), .D(\position1/n959 ), .Q(\position1/n1611 ) );
  NAND22 U2385 ( .A(\position1/x_sum [24]), .B(n673), .Q(\position1/n957 ) );
  NAND22 U2386 ( .A(\position1/N1201 ), .B(n636), .Q(\position1/n959 ) );
  AOI221 U2387 ( .A(\position1/N509 ), .B(n511), .C(\position1/N928 ), .D(n639), .Q(\position1/n958 ) );
  NOR31 U2388 ( .A(n1364), .B(n1363), .C(n1362), .Q(n1365) );
  NAND22 U2389 ( .A(\gensync1/N170 ), .B(\gensync1/N168 ), .Q(n1362) );
  NAND31 U2390 ( .A(\gensync1/N165 ), .B(\gensync1/N166 ), .C(\gensync1/N169 ), 
        .Q(n1363) );
  NAND41 U2391 ( .A(\gensync1/N173 ), .B(\gensync1/N171 ), .C(\gensync1/N172 ), 
        .D(\gensync1/N167 ), .Q(n1364) );
  NOR40 U2392 ( .A(n1369), .B(\gensync1/N166 ), .C(\gensync1/comptY[9] ), .D(
        \gensync1/N165 ), .Q(\gensync1/N132 ) );
  NOR21 U2393 ( .A(\gensync1/N167 ), .B(\gensync1/N168 ), .Q(n1366) );
  NAND22 U2394 ( .A(\gensync1/N169 ), .B(\gensync1/N170 ), .Q(n1367) );
  INV3 U2395 ( .A(\gensync1/n98 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [2]) );
  NAND22 U2396 ( .A(n814), .B(\gensync1/N138 ), .Q(\gensync1/n98 ) );
  XOR21 U2397 ( .A(\gensync1/N173 ), .B(\gensync1/N172 ), .Q(\gensync1/N138 )
         );
  NAND31 U2398 ( .A(\gensync1/N172 ), .B(\gensync1/N173 ), .C(\gensync1/N171 ), 
        .Q(n1368) );
  NOR21 U2399 ( .A(n198), .B(n75), .Q(\position1/r409/carry [13]) );
  INV3 U2400 ( .A(\position1/r409/carry [12]), .Q(n198) );
  NOR21 U2401 ( .A(n182), .B(n81), .Q(\position1/r406/carry [13]) );
  INV3 U2402 ( .A(\position1/r406/carry [12]), .Q(n182) );
  NOR21 U2403 ( .A(n196), .B(n68), .Q(\position1/r409/carry [11]) );
  INV3 U2404 ( .A(\position1/r409/carry [10]), .Q(n196) );
  NOR21 U2405 ( .A(n180), .B(n69), .Q(\position1/r406/carry [11]) );
  INV3 U2406 ( .A(\position1/r406/carry [10]), .Q(n180) );
  NOR21 U2407 ( .A(n195), .B(n50), .Q(\position1/r409/carry [10]) );
  INV3 U2408 ( .A(\position1/r409/carry [9]), .Q(n195) );
  NOR21 U2409 ( .A(n179), .B(n51), .Q(\position1/r406/carry [10]) );
  INV3 U2410 ( .A(\position1/r406/carry [9]), .Q(n179) );
  NOR21 U2411 ( .A(n197), .B(n58), .Q(\position1/r409/carry [12]) );
  INV3 U2412 ( .A(\position1/r409/carry [11]), .Q(n197) );
  NOR21 U2413 ( .A(n181), .B(n65), .Q(\position1/r406/carry [12]) );
  INV3 U2414 ( .A(\position1/r406/carry [11]), .Q(n181) );
  INV3 U2415 ( .A(\gensync1/N66 ), .Q(n872) );
  NOR40 U2416 ( .A(\gensync1/N174 ), .B(\gensync1/N175 ), .C(\gensync1/N176 ), 
        .D(n1383), .Q(\gensync1/N66 ) );
  NOR21 U2417 ( .A(n1382), .B(n6), .Q(n1383) );
  AOI311 U2418 ( .A(\gensync1/N180 ), .B(\gensync1/N181 ), .C(\gensync1/N179 ), 
        .D(\gensync1/N178 ), .Q(n1382) );
  AOI221 U2419 ( .A(\position1/N428 ), .B(n644), .C(\position1/N655 ), .D(n647), .Q(\position1/n860 ) );
  XOR21 U2420 ( .A(\position1/y_sum [23]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [23]), .Q(\position1/N655 )
         );
  XOR21 U2421 ( .A(\position1/N378 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [23]), .Q(
        \position1/N428 ) );
  AOI221 U2422 ( .A(\position1/N353 ), .B(n642), .C(\position1/N630 ), .D(n646), .Q(\position1/n960 ) );
  XOR21 U2423 ( .A(\position1/x_sum [23]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [23]), .Q(\position1/N630 )
         );
  XOR21 U2424 ( .A(\position1/N303 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [23]), .Q(
        \position1/N353 ) );
  AOI221 U2425 ( .A(\position1/N352 ), .B(n642), .C(\position1/N629 ), .D(n646), .Q(\position1/n964 ) );
  XOR21 U2426 ( .A(\position1/x_sum [22]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [22]), .Q(\position1/N629 )
         );
  XOR21 U2427 ( .A(\position1/N302 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [22]), .Q(
        \position1/N352 ) );
  AOI221 U2428 ( .A(\position1/N429 ), .B(n644), .C(\position1/N656 ), .D(n647), .Q(\position1/n852 ) );
  XOR21 U2429 ( .A(\position1/dp_cluster_5/add_179_aco/carry [24]), .B(
        \position1/y_sum [24]), .Q(\position1/N656 ) );
  XOR21 U2430 ( .A(\position1/dp_cluster_6/add_0_root_add_171_3/carry [24]), 
        .B(\position1/N379 ), .Q(\position1/N429 ) );
  NOR21 U2431 ( .A(n410), .B(n52), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [24]) );
  AOI221 U2432 ( .A(\position1/N354 ), .B(n642), .C(\position1/N631 ), .D(n646), .Q(\position1/n956 ) );
  XOR21 U2433 ( .A(\position1/dp_cluster_4/add_178_aco/carry [24]), .B(
        \position1/x_sum [24]), .Q(\position1/N631 ) );
  XOR21 U2434 ( .A(\position1/dp_cluster_7/add_0_root_add_170_3/carry [24]), 
        .B(\position1/N304 ), .Q(\position1/N354 ) );
  NOR21 U2435 ( .A(n395), .B(n59), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [24]) );
  INV3 U2436 ( .A(\gensync1/n105 ), .Q(n814) );
  NAND22 U2437 ( .A(\gensync1/n106 ), .B(\gensync1/N135 ), .Q(\gensync1/n105 )
         );
  NOR21 U2438 ( .A(\gensync1/comptY[9] ), .B(n1365), .Q(\gensync1/N135 ) );
  NOR21 U2439 ( .A(\gensync1/N132 ), .B(\gensync1/N129 ), .Q(\gensync1/n106 )
         );
  NOR21 U2440 ( .A(n505), .B(n10), .Q(n2133) );
  NOR21 U2441 ( .A(n505), .B(n1), .Q(n2134) );
  NOR21 U2442 ( .A(n194), .B(n96), .Q(\position1/r409/carry [1]) );
  INV3 U2443 ( .A(cam_y[0]), .Q(n194) );
  AOI2111 U2444 ( .A(\gensync1/N176 ), .B(n870), .C(\gensync1/N174 ), .D(
        \gensync1/N175 ), .Q(\gensync1/N69 ) );
  INV3 U2445 ( .A(n1381), .Q(n870) );
  NOR40 U2446 ( .A(\gensync1/N177 ), .B(\gensync1/N178 ), .C(\gensync1/N179 ), 
        .D(n871), .Q(n1381) );
  INV3 U2447 ( .A(n1380), .Q(n871) );
  NOR21 U2448 ( .A(n199), .B(n57), .Q(\position1/r409/carry [14]) );
  INV3 U2449 ( .A(\position1/r409/carry [13]), .Q(n199) );
  NOR21 U2450 ( .A(n183), .B(n64), .Q(\position1/r406/carry [14]) );
  INV3 U2451 ( .A(\position1/r406/carry [13]), .Q(n183) );
  NOR21 U2452 ( .A(n201), .B(n56), .Q(\position1/r409/carry [16]) );
  INV3 U2453 ( .A(\position1/r409/carry [15]), .Q(n201) );
  NOR21 U2454 ( .A(n185), .B(n63), .Q(\position1/r406/carry [16]) );
  INV3 U2455 ( .A(\position1/r406/carry [15]), .Q(n185) );
  NOR21 U2456 ( .A(n203), .B(n55), .Q(\position1/r409/carry [18]) );
  INV3 U2457 ( .A(\position1/r409/carry [17]), .Q(n203) );
  NOR21 U2458 ( .A(n187), .B(n62), .Q(\position1/r406/carry [18]) );
  INV3 U2459 ( .A(\position1/r406/carry [17]), .Q(n187) );
  NOR21 U2460 ( .A(n205), .B(n54), .Q(\position1/r409/carry [20]) );
  INV3 U2461 ( .A(\position1/r409/carry [19]), .Q(n205) );
  NOR21 U2462 ( .A(n189), .B(n61), .Q(\position1/r406/carry [20]) );
  INV3 U2463 ( .A(\position1/r406/carry [19]), .Q(n189) );
  NOR21 U2464 ( .A(n207), .B(n53), .Q(\position1/r409/carry [22]) );
  INV3 U2465 ( .A(\position1/r409/carry [21]), .Q(n207) );
  NOR21 U2466 ( .A(n191), .B(n60), .Q(\position1/r406/carry [22]) );
  INV3 U2467 ( .A(\position1/r406/carry [21]), .Q(n191) );
  XOR21 U2468 ( .A(\position1/r406/carry [24]), .B(\position1/x_sum [24]), .Q(
        \position1/N304 ) );
  NOR21 U2469 ( .A(n193), .B(n59), .Q(\position1/r406/carry [24]) );
  INV3 U2470 ( .A(\position1/r406/carry [23]), .Q(n193) );
  NOR21 U2471 ( .A(n178), .B(n97), .Q(\position1/r406/carry [1]) );
  INV3 U2472 ( .A(n503), .Q(n178) );
  NOR21 U2473 ( .A(n200), .B(n74), .Q(\position1/r409/carry [15]) );
  INV3 U2474 ( .A(\position1/r409/carry [14]), .Q(n200) );
  NOR21 U2475 ( .A(n184), .B(n80), .Q(\position1/r406/carry [15]) );
  INV3 U2476 ( .A(\position1/r406/carry [14]), .Q(n184) );
  NOR21 U2477 ( .A(n202), .B(n73), .Q(\position1/r409/carry [17]) );
  INV3 U2478 ( .A(\position1/r409/carry [16]), .Q(n202) );
  NOR21 U2479 ( .A(n186), .B(n79), .Q(\position1/r406/carry [17]) );
  INV3 U2480 ( .A(\position1/r406/carry [16]), .Q(n186) );
  NOR21 U2481 ( .A(n204), .B(n72), .Q(\position1/r409/carry [19]) );
  INV3 U2482 ( .A(\position1/r409/carry [18]), .Q(n204) );
  NOR21 U2483 ( .A(n188), .B(n78), .Q(\position1/r406/carry [19]) );
  INV3 U2484 ( .A(\position1/r406/carry [18]), .Q(n188) );
  NOR21 U2485 ( .A(n206), .B(n71), .Q(\position1/r409/carry [21]) );
  INV3 U2486 ( .A(\position1/r409/carry [20]), .Q(n206) );
  NOR21 U2487 ( .A(n190), .B(n77), .Q(\position1/r406/carry [21]) );
  INV3 U2488 ( .A(\position1/r406/carry [20]), .Q(n190) );
  NOR21 U2489 ( .A(n208), .B(n70), .Q(\position1/r409/carry [23]) );
  INV3 U2490 ( .A(\position1/r409/carry [22]), .Q(n208) );
  NOR21 U2491 ( .A(n192), .B(n76), .Q(\position1/r406/carry [23]) );
  INV3 U2492 ( .A(\position1/r406/carry [22]), .Q(n192) );
  XOR21 U2493 ( .A(\position1/N1938 ), .B(cam_y[0]), .Q(\position1/N355 ) );
  XOR21 U2494 ( .A(\position1/N1521 ), .B(n503), .Q(\position1/N280 ) );
  INV3 U2495 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[8] ), .Q(
        n777) );
  NAND22 U2496 ( .A(n1361), .B(\position1/dp_cluster_6/N389 ), .Q(
        \position1/dp_cluster_5/mult_add_179_aco/PROD_not[8] ) );
  INV3 U2497 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[8] ), .Q(
        n867) );
  NAND22 U2498 ( .A(n1361), .B(\position1/dp_cluster_7/N314 ), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[8] ) );
  INV3 U2499 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[8] ), .Q(
        n868) );
  NAND22 U2500 ( .A(n1360), .B(\position1/dp_cluster_7/N314 ), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[8] ) );
  NAND41 U2501 ( .A(\position1/n868 ), .B(\position1/n869 ), .C(
        \position1/n870 ), .D(\position1/n871 ), .Q(\position1/n1589 ) );
  NAND22 U2502 ( .A(\position1/y_sum [21]), .B(n509), .Q(\position1/n869 ) );
  NAND22 U2503 ( .A(\position1/N1223 ), .B(n637), .Q(\position1/n871 ) );
  AOI221 U2504 ( .A(\position1/N556 ), .B(n512), .C(\position1/N1000 ), .D(
        n641), .Q(\position1/n870 ) );
  NAND41 U2505 ( .A(\position1/n864 ), .B(\position1/n865 ), .C(
        \position1/n866 ), .D(\position1/n867 ), .Q(\position1/n1588 ) );
  NAND22 U2506 ( .A(\position1/y_sum [22]), .B(n509), .Q(\position1/n865 ) );
  NAND22 U2507 ( .A(\position1/N1224 ), .B(n637), .Q(\position1/n867 ) );
  AOI221 U2508 ( .A(\position1/N557 ), .B(n512), .C(\position1/N1001 ), .D(
        n641), .Q(\position1/n866 ) );
  NAND41 U2509 ( .A(\position1/n972 ), .B(\position1/n973 ), .C(
        \position1/n974 ), .D(\position1/n975 ), .Q(\position1/n1615 ) );
  NAND22 U2510 ( .A(\position1/x_sum [20]), .B(n508), .Q(\position1/n973 ) );
  NAND22 U2511 ( .A(\position1/N1197 ), .B(n635), .Q(\position1/n975 ) );
  AOI221 U2512 ( .A(\position1/N505 ), .B(n511), .C(\position1/N924 ), .D(n639), .Q(\position1/n974 ) );
  NAND41 U2513 ( .A(\position1/n968 ), .B(\position1/n969 ), .C(
        \position1/n970 ), .D(\position1/n971 ), .Q(\position1/n1614 ) );
  NAND22 U2514 ( .A(\position1/x_sum [21]), .B(n508), .Q(\position1/n969 ) );
  NAND22 U2515 ( .A(\position1/N1198 ), .B(n635), .Q(\position1/n971 ) );
  AOI221 U2516 ( .A(\position1/N506 ), .B(n511), .C(\position1/N925 ), .D(n639), .Q(\position1/n970 ) );
  INV3 U2517 ( .A(\gensync1/n97 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [3]) );
  NAND22 U2518 ( .A(n814), .B(\gensync1/N139 ), .Q(\gensync1/n97 ) );
  XOR21 U2519 ( .A(\gensync1/sub_95_2_cf/carry[2] ), .B(\gensync1/N171 ), .Q(
        \gensync1/N139 ) );
  NOR21 U2520 ( .A(n396), .B(n50), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [10]) );
  INV3 U2521 ( .A(\position1/dp_cluster_5/add_179_aco/carry [9]), .Q(n396) );
  NOR21 U2522 ( .A(n381), .B(n51), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [10]) );
  INV3 U2523 ( .A(\position1/dp_cluster_4/add_178_aco/carry [9]), .Q(n381) );
  NOR21 U2524 ( .A(n398), .B(n58), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [12]) );
  INV3 U2525 ( .A(\position1/dp_cluster_5/add_179_aco/carry [11]), .Q(n398) );
  NOR21 U2526 ( .A(n383), .B(n65), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [12]) );
  INV3 U2527 ( .A(\position1/dp_cluster_4/add_178_aco/carry [11]), .Q(n383) );
  NOR21 U2528 ( .A(n321), .B(n65), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [12]) );
  INV3 U2529 ( .A(\position1/dp_cluster_0/add_196_aco/carry [11]), .Q(n321) );
  NAND22 U2530 ( .A(\gensync1/N174 ), .B(\gensync1/N175 ), .Q(\gensync1/N85 )
         );
  INV3 U2531 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[5] ), .Q(
        n860) );
  NAND22 U2532 ( .A(cam_x[5]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[5] ) );
  INV3 U2533 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[1] ), .Q(
        n807) );
  NOR21 U2534 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[0] ), .B(
        n96), .Q(\position1/dp_cluster_5/add_179_aco/carry [1]) );
  NAND22 U2535 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[1] )
         );
  INV3 U2536 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[4] ), .Q(
        n795) );
  NAND22 U2537 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[4] )
         );
  INV3 U2538 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[5] ), .Q(
        n791) );
  NAND22 U2539 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[5] )
         );
  INV3 U2540 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[4] ), .Q(
        n858) );
  NAND22 U2541 ( .A(cam_x[4]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[4] ) );
  INV3 U2542 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[4] ), .Q(
        n859) );
  NAND22 U2543 ( .A(cam_x[4]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[4] ) );
  INV3 U2544 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[5] ), .Q(
        n861) );
  NAND22 U2545 ( .A(cam_x[5]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[5] ) );
  INV3 U2546 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[6] ), .Q(
        n787) );
  NAND22 U2547 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[6] )
         );
  INV3 U2548 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[6] ), .Q(
        n862) );
  NAND22 U2549 ( .A(cam_x[6]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[6] ) );
  INV3 U2550 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[2] ), .Q(
        n803) );
  NAND22 U2551 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[2] )
         );
  INV3 U2552 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[2] ), .Q(
        n855) );
  NAND22 U2553 ( .A(n499), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[2] ) );
  INV3 U2554 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[2] ), .Q(
        n854) );
  NAND22 U2555 ( .A(cam_x[2]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[2] ) );
  INV3 U2556 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[6] ), .Q(
        n863) );
  NAND22 U2557 ( .A(cam_x[6]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[6] ) );
  INV3 U2558 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[7] ), .Q(
        n783) );
  NAND22 U2559 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[7] )
         );
  INV3 U2560 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[7] ), .Q(
        n865) );
  NAND22 U2561 ( .A(cam_x[7]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[7] ) );
  INV3 U2562 ( .A(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[3] ), .Q(
        n799) );
  NAND22 U2563 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), 
        .B(n1361), .Q(\position1/dp_cluster_5/mult_add_179_aco/PROD_not[3] )
         );
  INV3 U2564 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[3] ), .Q(
        n857) );
  NAND22 U2565 ( .A(n497), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[3] ) );
  INV3 U2566 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[3] ), .Q(
        n856) );
  NAND22 U2567 ( .A(cam_x[3]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[3] ) );
  INV3 U2568 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[7] ), .Q(
        n866) );
  NAND22 U2569 ( .A(cam_x[7]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[7] ) );
  AOI221 U2570 ( .A(\position1/N426 ), .B(n644), .C(\position1/N653 ), .D(n647), .Q(\position1/n868 ) );
  XOR21 U2571 ( .A(\position1/y_sum [21]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [21]), .Q(\position1/N653 )
         );
  XOR21 U2572 ( .A(\position1/N376 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [21]), .Q(
        \position1/N426 ) );
  AOI221 U2573 ( .A(\position1/N427 ), .B(n644), .C(\position1/N654 ), .D(n647), .Q(\position1/n864 ) );
  XOR21 U2574 ( .A(\position1/y_sum [22]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [22]), .Q(\position1/N654 )
         );
  XOR21 U2575 ( .A(\position1/N377 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [22]), .Q(
        \position1/N427 ) );
  AOI221 U2576 ( .A(\position1/N350 ), .B(n642), .C(\position1/N627 ), .D(n646), .Q(\position1/n972 ) );
  XOR21 U2577 ( .A(\position1/x_sum [20]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [20]), .Q(\position1/N627 )
         );
  XOR21 U2578 ( .A(\position1/N300 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [20]), .Q(
        \position1/N350 ) );
  AOI221 U2579 ( .A(\position1/N351 ), .B(n642), .C(\position1/N628 ), .D(n646), .Q(\position1/n968 ) );
  XOR21 U2580 ( .A(\position1/x_sum [21]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [21]), .Q(\position1/N628 )
         );
  XOR21 U2581 ( .A(\position1/N301 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [21]), .Q(
        \position1/N351 ) );
  NOR21 U2582 ( .A(n505), .B(n4), .Q(n2132) );
  NOR21 U2583 ( .A(n505), .B(n12), .Q(n2131) );
  INV3 U2584 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[1] ), .Q(
        n835) );
  NOR21 U2585 ( .A(\position1/dp_cluster_0/mult_add_196_aco/PROD_not[0] ), .B(
        n97), .Q(\position1/dp_cluster_0/add_196_aco/carry [1]) );
  NAND22 U2586 ( .A(cam_x[1]), .B(n1360), .Q(
        \position1/dp_cluster_0/mult_add_196_aco/PROD_not[1] ) );
  INV3 U2587 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[1] ), .Q(
        n834) );
  NOR21 U2588 ( .A(\position1/dp_cluster_4/mult_add_178_aco/PROD_not[0] ), .B(
        n97), .Q(\position1/dp_cluster_4/add_178_aco/carry [1]) );
  NAND22 U2589 ( .A(cam_x[1]), .B(n1361), .Q(
        \position1/dp_cluster_4/mult_add_178_aco/PROD_not[1] ) );
  NOR21 U2590 ( .A(n319), .B(n51), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [10]) );
  INV3 U2591 ( .A(\position1/dp_cluster_0/add_196_aco/carry [9]), .Q(n319) );
  NOR21 U2592 ( .A(n400), .B(n57), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [14]) );
  INV3 U2593 ( .A(\position1/dp_cluster_5/add_179_aco/carry [13]), .Q(n400) );
  NOR21 U2594 ( .A(n385), .B(n64), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [14]) );
  INV3 U2595 ( .A(\position1/dp_cluster_4/add_178_aco/carry [13]), .Q(n385) );
  NOR21 U2596 ( .A(n323), .B(n64), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [14]) );
  INV3 U2597 ( .A(\position1/dp_cluster_0/add_196_aco/carry [13]), .Q(n323) );
  NOR21 U2598 ( .A(n402), .B(n56), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [16]) );
  INV3 U2599 ( .A(\position1/dp_cluster_5/add_179_aco/carry [15]), .Q(n402) );
  NOR21 U2600 ( .A(n387), .B(n63), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [16]) );
  INV3 U2601 ( .A(\position1/dp_cluster_4/add_178_aco/carry [15]), .Q(n387) );
  NOR21 U2602 ( .A(n325), .B(n63), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [16]) );
  INV3 U2603 ( .A(\position1/dp_cluster_0/add_196_aco/carry [15]), .Q(n325) );
  NOR21 U2604 ( .A(n404), .B(n55), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [18]) );
  INV3 U2605 ( .A(\position1/dp_cluster_5/add_179_aco/carry [17]), .Q(n404) );
  NOR21 U2606 ( .A(n389), .B(n62), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [18]) );
  INV3 U2607 ( .A(\position1/dp_cluster_4/add_178_aco/carry [17]), .Q(n389) );
  NOR21 U2608 ( .A(n327), .B(n62), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [18]) );
  INV3 U2609 ( .A(\position1/dp_cluster_0/add_196_aco/carry [17]), .Q(n327) );
  NOR21 U2610 ( .A(n406), .B(n54), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [20]) );
  INV3 U2611 ( .A(\position1/dp_cluster_5/add_179_aco/carry [19]), .Q(n406) );
  NOR21 U2612 ( .A(n391), .B(n61), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [20]) );
  INV3 U2613 ( .A(\position1/dp_cluster_4/add_178_aco/carry [19]), .Q(n391) );
  NOR21 U2614 ( .A(n329), .B(n61), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [20]) );
  INV3 U2615 ( .A(\position1/dp_cluster_0/add_196_aco/carry [19]), .Q(n329) );
  NOR21 U2616 ( .A(n408), .B(n53), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [22]) );
  INV3 U2617 ( .A(\position1/dp_cluster_5/add_179_aco/carry [21]), .Q(n408) );
  NOR21 U2618 ( .A(n393), .B(n60), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [22]) );
  INV3 U2619 ( .A(\position1/dp_cluster_4/add_178_aco/carry [21]), .Q(n393) );
  NOR21 U2620 ( .A(n331), .B(n60), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [22]) );
  INV3 U2621 ( .A(\position1/dp_cluster_0/add_196_aco/carry [21]), .Q(n331) );
  XOR21 U2622 ( .A(\position1/r409/carry [24]), .B(\position1/y_sum [24]), .Q(
        \position1/N379 ) );
  NOR21 U2623 ( .A(n209), .B(n52), .Q(\position1/r409/carry [24]) );
  INV3 U2624 ( .A(\position1/r409/carry [23]), .Q(n209) );
  XOR21 U2625 ( .A(\position1/dp_cluster_0/add_196_aco/carry [24]), .B(
        \position1/x_sum [24]), .Q(\position1/N1201 ) );
  NOR21 U2626 ( .A(n333), .B(n59), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [24]) );
  INV3 U2627 ( .A(\position1/dp_cluster_0/add_196_aco/carry [23]), .Q(n333) );
  NOR21 U2628 ( .A(n397), .B(n68), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [11]) );
  INV3 U2629 ( .A(\position1/dp_cluster_5/add_179_aco/carry [10]), .Q(n397) );
  NOR21 U2630 ( .A(n382), .B(n69), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [11]) );
  INV3 U2631 ( .A(\position1/dp_cluster_4/add_178_aco/carry [10]), .Q(n382) );
  NOR21 U2632 ( .A(n320), .B(n69), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [11]) );
  INV3 U2633 ( .A(\position1/dp_cluster_0/add_196_aco/carry [10]), .Q(n320) );
  NOR21 U2634 ( .A(n399), .B(n75), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [13]) );
  INV3 U2635 ( .A(\position1/dp_cluster_5/add_179_aco/carry [12]), .Q(n399) );
  NOR21 U2636 ( .A(n384), .B(n81), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [13]) );
  INV3 U2637 ( .A(\position1/dp_cluster_4/add_178_aco/carry [12]), .Q(n384) );
  NOR21 U2638 ( .A(n322), .B(n81), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [13]) );
  INV3 U2639 ( .A(\position1/dp_cluster_0/add_196_aco/carry [12]), .Q(n322) );
  NOR21 U2640 ( .A(n401), .B(n74), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [15]) );
  INV3 U2641 ( .A(\position1/dp_cluster_5/add_179_aco/carry [14]), .Q(n401) );
  NOR21 U2642 ( .A(n386), .B(n80), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [15]) );
  INV3 U2643 ( .A(\position1/dp_cluster_4/add_178_aco/carry [14]), .Q(n386) );
  NOR21 U2644 ( .A(n324), .B(n80), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [15]) );
  INV3 U2645 ( .A(\position1/dp_cluster_0/add_196_aco/carry [14]), .Q(n324) );
  NOR21 U2646 ( .A(n403), .B(n73), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [17]) );
  INV3 U2647 ( .A(\position1/dp_cluster_5/add_179_aco/carry [16]), .Q(n403) );
  NOR21 U2648 ( .A(n388), .B(n79), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [17]) );
  INV3 U2649 ( .A(\position1/dp_cluster_4/add_178_aco/carry [16]), .Q(n388) );
  NOR21 U2650 ( .A(n326), .B(n79), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [17]) );
  INV3 U2651 ( .A(\position1/dp_cluster_0/add_196_aco/carry [16]), .Q(n326) );
  NOR21 U2652 ( .A(n405), .B(n72), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [19]) );
  INV3 U2653 ( .A(\position1/dp_cluster_5/add_179_aco/carry [18]), .Q(n405) );
  NOR21 U2654 ( .A(n390), .B(n78), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [19]) );
  INV3 U2655 ( .A(\position1/dp_cluster_4/add_178_aco/carry [18]), .Q(n390) );
  NOR21 U2656 ( .A(n328), .B(n78), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [19]) );
  INV3 U2657 ( .A(\position1/dp_cluster_0/add_196_aco/carry [18]), .Q(n328) );
  NOR21 U2658 ( .A(n407), .B(n71), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [21]) );
  INV3 U2659 ( .A(\position1/dp_cluster_5/add_179_aco/carry [20]), .Q(n407) );
  NOR21 U2660 ( .A(n392), .B(n77), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [21]) );
  INV3 U2661 ( .A(\position1/dp_cluster_4/add_178_aco/carry [20]), .Q(n392) );
  NOR21 U2662 ( .A(n330), .B(n77), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [21]) );
  INV3 U2663 ( .A(\position1/dp_cluster_0/add_196_aco/carry [20]), .Q(n330) );
  NOR21 U2664 ( .A(n409), .B(n70), .Q(
        \position1/dp_cluster_5/add_179_aco/carry [23]) );
  INV3 U2665 ( .A(\position1/dp_cluster_5/add_179_aco/carry [22]), .Q(n409) );
  NOR21 U2666 ( .A(n394), .B(n76), .Q(
        \position1/dp_cluster_4/add_178_aco/carry [23]) );
  INV3 U2667 ( .A(\position1/dp_cluster_4/add_178_aco/carry [22]), .Q(n394) );
  NOR21 U2668 ( .A(n332), .B(n76), .Q(
        \position1/dp_cluster_0/add_196_aco/carry [23]) );
  INV3 U2669 ( .A(\position1/dp_cluster_0/add_196_aco/carry [22]), .Q(n332) );
  NAND31 U2670 ( .A(\position1/n1147 ), .B(\position1/n357 ), .C(
        \position1/n1187 ), .Q(\position1/n1145 ) );
  NAND31 U2671 ( .A(\position1/n1147 ), .B(\position1/gi [5]), .C(
        \position1/n1187 ), .Q(\position1/n1151 ) );
  NOR40 U2672 ( .A(\position1/n356 ), .B(\position1/n358 ), .C(
        \position1/gi [0]), .D(\position1/gi [2]), .Q(\position1/n1187 ) );
  INV3 U2673 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[8] ), .Q(
        n778) );
  NAND22 U2674 ( .A(n1360), .B(\position1/dp_cluster_6/N389 ), .Q(
        \position1/dp_cluster_1/mult_add_197_aco/PROD_not[8] ) );
  NAND41 U2675 ( .A(\position1/n880 ), .B(\position1/n881 ), .C(
        \position1/n882 ), .D(\position1/n883 ), .Q(\position1/n1592 ) );
  NAND22 U2676 ( .A(\position1/y_sum [18]), .B(n509), .Q(\position1/n881 ) );
  NAND22 U2677 ( .A(\position1/N1220 ), .B(n637), .Q(\position1/n883 ) );
  AOI221 U2678 ( .A(\position1/N553 ), .B(n512), .C(\position1/N997 ), .D(n641), .Q(\position1/n882 ) );
  NAND41 U2679 ( .A(\position1/n876 ), .B(\position1/n877 ), .C(
        \position1/n878 ), .D(\position1/n879 ), .Q(\position1/n1591 ) );
  NAND22 U2680 ( .A(\position1/y_sum [19]), .B(n509), .Q(\position1/n877 ) );
  NAND22 U2681 ( .A(\position1/N1221 ), .B(n637), .Q(\position1/n879 ) );
  AOI221 U2682 ( .A(\position1/N554 ), .B(n512), .C(\position1/N998 ), .D(n641), .Q(\position1/n878 ) );
  NAND41 U2683 ( .A(\position1/n872 ), .B(\position1/n873 ), .C(
        \position1/n874 ), .D(\position1/n875 ), .Q(\position1/n1590 ) );
  NAND22 U2684 ( .A(\position1/y_sum [20]), .B(n509), .Q(\position1/n873 ) );
  NAND22 U2685 ( .A(\position1/N1222 ), .B(n637), .Q(\position1/n875 ) );
  AOI221 U2686 ( .A(\position1/N555 ), .B(n512), .C(\position1/N999 ), .D(n641), .Q(\position1/n874 ) );
  NAND41 U2687 ( .A(\position1/n980 ), .B(\position1/n981 ), .C(
        \position1/n982 ), .D(\position1/n983 ), .Q(\position1/n1617 ) );
  NAND22 U2688 ( .A(\position1/x_sum [18]), .B(n508), .Q(\position1/n981 ) );
  NAND22 U2689 ( .A(\position1/N1195 ), .B(n635), .Q(\position1/n983 ) );
  AOI221 U2690 ( .A(\position1/N503 ), .B(n511), .C(\position1/N922 ), .D(n639), .Q(\position1/n982 ) );
  NAND41 U2691 ( .A(\position1/n976 ), .B(\position1/n977 ), .C(
        \position1/n978 ), .D(\position1/n979 ), .Q(\position1/n1616 ) );
  NAND22 U2692 ( .A(\position1/x_sum [19]), .B(n508), .Q(\position1/n977 ) );
  NAND22 U2693 ( .A(\position1/N1196 ), .B(n635), .Q(\position1/n979 ) );
  AOI221 U2694 ( .A(\position1/N504 ), .B(n511), .C(\position1/N923 ), .D(n639), .Q(\position1/n978 ) );
  INV3 U2695 ( .A(\gensync1/n96 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [4]) );
  NAND22 U2696 ( .A(n814), .B(\gensync1/N140 ), .Q(\gensync1/n96 ) );
  XOR21 U2697 ( .A(\gensync1/sub_95_2_cf/carry[3] ), .B(\gensync1/N170 ), .Q(
        \gensync1/N140 ) );
  INV3 U2698 ( .A(\gensync1/n95 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [5]) );
  NAND22 U2699 ( .A(n814), .B(\gensync1/N141 ), .Q(\gensync1/n95 ) );
  XOR21 U2700 ( .A(\gensync1/sub_95_2_cf/carry[4] ), .B(\gensync1/N169 ), .Q(
        \gensync1/N141 ) );
  NOR21 U2701 ( .A(n336), .B(n58), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [12]) );
  INV3 U2702 ( .A(\position1/dp_cluster_1/add_197_aco/carry [11]), .Q(n336) );
  NOR21 U2703 ( .A(n9), .B(n3), .Q(\gensync1/sub_95_2_cf/carry[2] ) );
  NOR21 U2704 ( .A(n8), .B(n463), .Q(\gensync1/sub_95_2_cf/carry[3] ) );
  INV3 U2705 ( .A(\gensync1/sub_95_2_cf/carry[2] ), .Q(n463) );
  XOR21 U2706 ( .A(\position1/y_sum [22]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [22]), .Q(\position1/N1224 )
         );
  XOR21 U2707 ( .A(\position1/x_sum [22]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [22]), .Q(\position1/N1199 )
         );
  XOR21 U2708 ( .A(\position1/y_sum [23]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [23]), .Q(\position1/N1225 )
         );
  XOR21 U2709 ( .A(\position1/x_sum [23]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [23]), .Q(\position1/N1200 )
         );
  INV3 U2710 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[1] ), .Q(
        n808) );
  NOR21 U2711 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[0] ), .B(
        n96), .Q(\position1/dp_cluster_1/add_197_aco/carry [1]) );
  NAND22 U2712 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[1] )
         );
  INV3 U2713 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[4] ), .Q(
        n796) );
  NAND22 U2714 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [5]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[4] )
         );
  INV3 U2715 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[5] ), .Q(
        n792) );
  NAND22 U2716 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [6]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[5] )
         );
  INV3 U2717 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[2] ), .Q(
        n804) );
  NAND22 U2718 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [3]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[2] )
         );
  INV3 U2719 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[6] ), .Q(
        n788) );
  NAND22 U2720 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [7]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[6] )
         );
  INV3 U2721 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[3] ), .Q(
        n800) );
  NAND22 U2722 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[3] )
         );
  INV3 U2723 ( .A(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[7] ), .Q(
        n784) );
  NAND22 U2724 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [8]), 
        .B(n1360), .Q(\position1/dp_cluster_1/mult_add_197_aco/PROD_not[7] )
         );
  AOI221 U2725 ( .A(\position1/N423 ), .B(n644), .C(\position1/N650 ), .D(n647), .Q(\position1/n880 ) );
  XOR21 U2726 ( .A(\position1/y_sum [18]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [18]), .Q(\position1/N650 )
         );
  XOR21 U2727 ( .A(\position1/N373 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [18]), .Q(
        \position1/N423 ) );
  AOI221 U2728 ( .A(\position1/N424 ), .B(n644), .C(\position1/N651 ), .D(n647), .Q(\position1/n876 ) );
  XOR21 U2729 ( .A(\position1/y_sum [19]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [19]), .Q(\position1/N651 )
         );
  XOR21 U2730 ( .A(\position1/N374 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [19]), .Q(
        \position1/N424 ) );
  AOI221 U2731 ( .A(\position1/N425 ), .B(n644), .C(\position1/N652 ), .D(n647), .Q(\position1/n872 ) );
  XOR21 U2732 ( .A(\position1/y_sum [20]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [20]), .Q(\position1/N652 )
         );
  XOR21 U2733 ( .A(\position1/N375 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [20]), .Q(
        \position1/N425 ) );
  AOI221 U2734 ( .A(\position1/N348 ), .B(n642), .C(\position1/N625 ), .D(n646), .Q(\position1/n980 ) );
  XOR21 U2735 ( .A(\position1/x_sum [18]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [18]), .Q(\position1/N625 )
         );
  XOR21 U2736 ( .A(\position1/N298 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [18]), .Q(
        \position1/N348 ) );
  AOI221 U2737 ( .A(\position1/N349 ), .B(n642), .C(\position1/N626 ), .D(n646), .Q(\position1/n976 ) );
  XOR21 U2738 ( .A(\position1/x_sum [19]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [19]), .Q(\position1/N626 )
         );
  XOR21 U2739 ( .A(\position1/N299 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [19]), .Q(
        \position1/N349 ) );
  NOR21 U2740 ( .A(n334), .B(n50), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [10]) );
  INV3 U2741 ( .A(\position1/dp_cluster_1/add_197_aco/carry [9]), .Q(n334) );
  NOR21 U2742 ( .A(n338), .B(n57), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [14]) );
  INV3 U2743 ( .A(\position1/dp_cluster_1/add_197_aco/carry [13]), .Q(n338) );
  NOR21 U2744 ( .A(n340), .B(n56), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [16]) );
  INV3 U2745 ( .A(\position1/dp_cluster_1/add_197_aco/carry [15]), .Q(n340) );
  NOR21 U2746 ( .A(n342), .B(n55), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [18]) );
  INV3 U2747 ( .A(\position1/dp_cluster_1/add_197_aco/carry [17]), .Q(n342) );
  NOR21 U2748 ( .A(n344), .B(n54), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [20]) );
  INV3 U2749 ( .A(\position1/dp_cluster_1/add_197_aco/carry [19]), .Q(n344) );
  NOR21 U2750 ( .A(n346), .B(n53), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [22]) );
  INV3 U2751 ( .A(\position1/dp_cluster_1/add_197_aco/carry [21]), .Q(n346) );
  XOR21 U2752 ( .A(\position1/dp_cluster_1/add_197_aco/carry [24]), .B(
        \position1/y_sum [24]), .Q(\position1/N1226 ) );
  NOR21 U2753 ( .A(n348), .B(n52), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [24]) );
  INV3 U2754 ( .A(\position1/dp_cluster_1/add_197_aco/carry [23]), .Q(n348) );
  NOR21 U2755 ( .A(n335), .B(n68), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [11]) );
  INV3 U2756 ( .A(\position1/dp_cluster_1/add_197_aco/carry [10]), .Q(n335) );
  NOR21 U2757 ( .A(n337), .B(n75), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [13]) );
  INV3 U2758 ( .A(\position1/dp_cluster_1/add_197_aco/carry [12]), .Q(n337) );
  NOR21 U2759 ( .A(n339), .B(n74), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [15]) );
  INV3 U2760 ( .A(\position1/dp_cluster_1/add_197_aco/carry [14]), .Q(n339) );
  NOR21 U2761 ( .A(n341), .B(n73), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [17]) );
  INV3 U2762 ( .A(\position1/dp_cluster_1/add_197_aco/carry [16]), .Q(n341) );
  NOR21 U2763 ( .A(n343), .B(n72), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [19]) );
  INV3 U2764 ( .A(\position1/dp_cluster_1/add_197_aco/carry [18]), .Q(n343) );
  NOR21 U2765 ( .A(n345), .B(n71), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [21]) );
  INV3 U2766 ( .A(\position1/dp_cluster_1/add_197_aco/carry [20]), .Q(n345) );
  NOR21 U2767 ( .A(n347), .B(n70), .Q(
        \position1/dp_cluster_1/add_197_aco/carry [23]) );
  INV3 U2768 ( .A(\position1/dp_cluster_1/add_197_aco/carry [22]), .Q(n347) );
  NOR31 U2769 ( .A(\position1/gi [3]), .B(\position1/gi [7]), .C(
        \position1/gi [1]), .Q(\position1/n1147 ) );
  NAND41 U2770 ( .A(\position1/n888 ), .B(\position1/n889 ), .C(
        \position1/n890 ), .D(\position1/n891 ), .Q(\position1/n1594 ) );
  NAND22 U2771 ( .A(\position1/y_sum [16]), .B(n509), .Q(\position1/n889 ) );
  NAND22 U2772 ( .A(\position1/N1218 ), .B(n637), .Q(\position1/n891 ) );
  AOI221 U2773 ( .A(\position1/N551 ), .B(n512), .C(\position1/N995 ), .D(n641), .Q(\position1/n890 ) );
  NAND41 U2774 ( .A(\position1/n884 ), .B(\position1/n885 ), .C(
        \position1/n886 ), .D(\position1/n887 ), .Q(\position1/n1593 ) );
  NAND22 U2775 ( .A(\position1/y_sum [17]), .B(n509), .Q(\position1/n885 ) );
  NAND22 U2776 ( .A(\position1/N1219 ), .B(n637), .Q(\position1/n887 ) );
  AOI221 U2777 ( .A(\position1/N552 ), .B(n512), .C(\position1/N996 ), .D(n641), .Q(\position1/n886 ) );
  NAND41 U2778 ( .A(\position1/n988 ), .B(\position1/n989 ), .C(
        \position1/n990 ), .D(\position1/n991 ), .Q(\position1/n1619 ) );
  NAND22 U2779 ( .A(\position1/x_sum [16]), .B(n508), .Q(\position1/n989 ) );
  NAND22 U2780 ( .A(\position1/N1193 ), .B(n635), .Q(\position1/n991 ) );
  AOI221 U2781 ( .A(\position1/N501 ), .B(n511), .C(\position1/N920 ), .D(n639), .Q(\position1/n990 ) );
  NAND41 U2782 ( .A(\position1/n984 ), .B(\position1/n985 ), .C(
        \position1/n986 ), .D(\position1/n987 ), .Q(\position1/n1618 ) );
  NAND22 U2783 ( .A(\position1/x_sum [17]), .B(n508), .Q(\position1/n985 ) );
  NAND22 U2784 ( .A(\position1/N1194 ), .B(n635), .Q(\position1/n987 ) );
  AOI221 U2785 ( .A(\position1/N502 ), .B(n511), .C(\position1/N921 ), .D(n639), .Q(\position1/n986 ) );
  INV3 U2786 ( .A(\gensync1/n93 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [7]) );
  NAND22 U2787 ( .A(n814), .B(\gensync1/N143 ), .Q(\gensync1/n93 ) );
  XNR21 U2788 ( .A(\gensync1/sub_95_2_cf/carry[6] ), .B(\gensync1/N167 ), .Q(
        \gensync1/N143 ) );
  INV3 U2789 ( .A(\gensync1/n92 ), .Q(
        \position1/dp_cluster_6/add_1_root_add_171_3/carry [8]) );
  NAND22 U2790 ( .A(n814), .B(\gensync1/N144 ), .Q(\gensync1/n92 ) );
  XNR21 U2791 ( .A(\gensync1/sub_95_2_cf/carry[7] ), .B(\gensync1/N166 ), .Q(
        \gensync1/N144 ) );
  NAND22 U2792 ( .A(n814), .B(\gensync1/N142 ), .Q(\gensync1/n94 ) );
  XNR21 U2793 ( .A(\gensync1/sub_95_2_cf/carry[5] ), .B(\gensync1/N168 ), .Q(
        \gensync1/N142 ) );
  NOR21 U2794 ( .A(n11), .B(n464), .Q(\gensync1/sub_95_2_cf/carry[4] ) );
  INV3 U2795 ( .A(\gensync1/sub_95_2_cf/carry[3] ), .Q(n464) );
  XOR21 U2796 ( .A(\position1/y_sum [20]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [20]), .Q(\position1/N1222 )
         );
  XOR21 U2797 ( .A(\position1/x_sum [20]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [20]), .Q(\position1/N1197 )
         );
  XOR21 U2798 ( .A(\position1/y_sum [21]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [21]), .Q(\position1/N1223 )
         );
  XOR21 U2799 ( .A(\position1/x_sum [19]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [19]), .Q(\position1/N1196 )
         );
  XOR21 U2800 ( .A(\position1/x_sum [21]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [21]), .Q(\position1/N1198 )
         );
  AOI221 U2801 ( .A(\position1/N421 ), .B(n644), .C(\position1/N648 ), .D(n647), .Q(\position1/n888 ) );
  XOR21 U2802 ( .A(\position1/y_sum [16]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [16]), .Q(\position1/N648 )
         );
  XOR21 U2803 ( .A(\position1/N371 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [16]), .Q(
        \position1/N421 ) );
  AOI221 U2804 ( .A(\position1/N422 ), .B(n644), .C(\position1/N649 ), .D(n647), .Q(\position1/n884 ) );
  XOR21 U2805 ( .A(\position1/y_sum [17]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [17]), .Q(\position1/N649 )
         );
  XOR21 U2806 ( .A(\position1/N372 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [17]), .Q(
        \position1/N422 ) );
  AOI221 U2807 ( .A(\position1/N346 ), .B(n642), .C(\position1/N623 ), .D(n646), .Q(\position1/n988 ) );
  XOR21 U2808 ( .A(\position1/x_sum [16]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [16]), .Q(\position1/N623 )
         );
  XOR21 U2809 ( .A(\position1/N296 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [16]), .Q(
        \position1/N346 ) );
  AOI221 U2810 ( .A(\position1/N347 ), .B(n642), .C(\position1/N624 ), .D(n646), .Q(\position1/n984 ) );
  XOR21 U2811 ( .A(\position1/x_sum [17]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [17]), .Q(\position1/N624 )
         );
  XOR21 U2812 ( .A(\position1/N297 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [17]), .Q(
        \position1/N347 ) );
  NOR21 U2813 ( .A(n505), .B(n14), .Q(n2129) );
  INV3 U2814 ( .A(n161), .Q(\gensync1/sub_95_2_cf/carry[6] ) );
  NOR21 U2815 ( .A(\gensync1/N168 ), .B(\gensync1/sub_95_2_cf/carry[5] ), .Q(
        n161) );
  INV3 U2816 ( .A(n162), .Q(\gensync1/sub_95_2_cf/carry[7] ) );
  NOR21 U2817 ( .A(\gensync1/N167 ), .B(\gensync1/sub_95_2_cf/carry[6] ), .Q(
        n162) );
  NOR21 U2818 ( .A(n13), .B(n465), .Q(\gensync1/sub_95_2_cf/carry[5] ) );
  INV3 U2819 ( .A(\gensync1/sub_95_2_cf/carry[4] ), .Q(n465) );
  NAND41 U2820 ( .A(\position1/n896 ), .B(\position1/n897 ), .C(
        \position1/n898 ), .D(\position1/n899 ), .Q(\position1/n1596 ) );
  NAND22 U2821 ( .A(\position1/y_sum [14]), .B(n509), .Q(\position1/n897 ) );
  NAND22 U2822 ( .A(\position1/N1216 ), .B(n637), .Q(\position1/n899 ) );
  AOI221 U2823 ( .A(\position1/N549 ), .B(n512), .C(\position1/N993 ), .D(n641), .Q(\position1/n898 ) );
  NAND41 U2824 ( .A(\position1/n892 ), .B(\position1/n893 ), .C(
        \position1/n894 ), .D(\position1/n895 ), .Q(\position1/n1595 ) );
  NAND22 U2825 ( .A(\position1/y_sum [15]), .B(n509), .Q(\position1/n893 ) );
  NAND22 U2826 ( .A(\position1/N1217 ), .B(n637), .Q(\position1/n895 ) );
  AOI221 U2827 ( .A(\position1/N550 ), .B(n512), .C(\position1/N994 ), .D(n641), .Q(\position1/n894 ) );
  NAND41 U2828 ( .A(\position1/n1000 ), .B(\position1/n1001 ), .C(
        \position1/n1002 ), .D(\position1/n1003 ), .Q(\position1/n1622 ) );
  NAND22 U2829 ( .A(\position1/x_sum [13]), .B(n508), .Q(\position1/n1001 ) );
  NAND22 U2830 ( .A(\position1/N1190 ), .B(n635), .Q(\position1/n1003 ) );
  AOI221 U2831 ( .A(\position1/N498 ), .B(n511), .C(\position1/N917 ), .D(n639), .Q(\position1/n1002 ) );
  NAND41 U2832 ( .A(\position1/n996 ), .B(\position1/n997 ), .C(
        \position1/n998 ), .D(\position1/n999 ), .Q(\position1/n1621 ) );
  NAND22 U2833 ( .A(\position1/x_sum [14]), .B(n508), .Q(\position1/n997 ) );
  NAND22 U2834 ( .A(\position1/N1191 ), .B(n635), .Q(\position1/n999 ) );
  AOI221 U2835 ( .A(\position1/N499 ), .B(n511), .C(\position1/N918 ), .D(n639), .Q(\position1/n998 ) );
  NAND41 U2836 ( .A(\position1/n992 ), .B(\position1/n993 ), .C(
        \position1/n994 ), .D(\position1/n995 ), .Q(\position1/n1620 ) );
  NAND22 U2837 ( .A(\position1/x_sum [15]), .B(n508), .Q(\position1/n993 ) );
  NAND22 U2838 ( .A(\position1/N1192 ), .B(n635), .Q(\position1/n995 ) );
  AOI221 U2839 ( .A(\position1/N500 ), .B(n511), .C(\position1/N919 ), .D(n639), .Q(\position1/n994 ) );
  NOR21 U2840 ( .A(\gensync1/N166 ), .B(\gensync1/sub_95_2_cf/carry[7] ), .Q(
        n163) );
  AOI221 U2841 ( .A(\position1/N344 ), .B(n642), .C(\position1/N621 ), .D(n646), .Q(\position1/n996 ) );
  XOR21 U2842 ( .A(\position1/x_sum [14]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [14]), .Q(\position1/N621 )
         );
  XOR21 U2843 ( .A(\position1/N294 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [14]), .Q(
        \position1/N344 ) );
  INV3 U2844 ( .A(\gensync1/n91 ), .Q(\position1/dp_cluster_6/N389 ) );
  NAND22 U2845 ( .A(n814), .B(\gensync1/N145 ), .Q(\gensync1/n91 ) );
  XNR21 U2846 ( .A(\gensync1/N165 ), .B(\gensync1/sub_95_2_cf/carry[8] ), .Q(
        \gensync1/N145 ) );
  INV3 U2847 ( .A(n163), .Q(\gensync1/sub_95_2_cf/carry[8] ) );
  XOR21 U2848 ( .A(\position1/y_sum [18]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [18]), .Q(\position1/N1220 )
         );
  XOR21 U2849 ( .A(\position1/x_sum [18]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [18]), .Q(\position1/N1195 )
         );
  XOR21 U2850 ( .A(\position1/y_sum [19]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [19]), .Q(\position1/N1221 )
         );
  XOR21 U2851 ( .A(\position1/x_sum [17]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [17]), .Q(\position1/N1194 )
         );
  AOI221 U2852 ( .A(\position1/N419 ), .B(n644), .C(\position1/N646 ), .D(n647), .Q(\position1/n896 ) );
  XOR21 U2853 ( .A(\position1/y_sum [14]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [14]), .Q(\position1/N646 )
         );
  XOR21 U2854 ( .A(\position1/N369 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [14]), .Q(
        \position1/N419 ) );
  AOI221 U2855 ( .A(\position1/N420 ), .B(n644), .C(\position1/N647 ), .D(n647), .Q(\position1/n892 ) );
  XOR21 U2856 ( .A(\position1/y_sum [15]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [15]), .Q(\position1/N647 )
         );
  XOR21 U2857 ( .A(\position1/N370 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [15]), .Q(
        \position1/N420 ) );
  AOI221 U2858 ( .A(\position1/N343 ), .B(n642), .C(\position1/N620 ), .D(n646), .Q(\position1/n1000 ) );
  XOR21 U2859 ( .A(\position1/x_sum [13]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [13]), .Q(\position1/N620 )
         );
  XOR21 U2860 ( .A(\position1/N293 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [13]), .Q(
        \position1/N343 ) );
  AOI221 U2861 ( .A(\position1/N345 ), .B(n642), .C(\position1/N622 ), .D(n646), .Q(\position1/n992 ) );
  XOR21 U2862 ( .A(\position1/x_sum [15]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [15]), .Q(\position1/N622 )
         );
  XOR21 U2863 ( .A(\position1/N295 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [15]), .Q(
        \position1/N345 ) );
  NOR21 U2864 ( .A(n505), .B(n15), .Q(n2127) );
  NAND41 U2865 ( .A(\position1/n904 ), .B(\position1/n905 ), .C(
        \position1/n906 ), .D(\position1/n907 ), .Q(\position1/n1598 ) );
  NAND22 U2866 ( .A(\position1/y_sum [12]), .B(n509), .Q(\position1/n905 ) );
  NAND22 U2867 ( .A(\position1/N1214 ), .B(n637), .Q(\position1/n907 ) );
  AOI221 U2868 ( .A(\position1/N547 ), .B(n740), .C(\position1/N991 ), .D(n640), .Q(\position1/n906 ) );
  NAND41 U2869 ( .A(\position1/n900 ), .B(\position1/n901 ), .C(
        \position1/n902 ), .D(\position1/n903 ), .Q(\position1/n1597 ) );
  NAND22 U2870 ( .A(\position1/y_sum [13]), .B(n509), .Q(\position1/n901 ) );
  NAND22 U2871 ( .A(\position1/N1215 ), .B(n637), .Q(\position1/n903 ) );
  AOI221 U2872 ( .A(\position1/N548 ), .B(n740), .C(\position1/N992 ), .D(n640), .Q(\position1/n902 ) );
  NAND41 U2873 ( .A(\position1/n1008 ), .B(\position1/n1009 ), .C(
        \position1/n1010 ), .D(\position1/n1011 ), .Q(\position1/n1624 ) );
  NAND22 U2874 ( .A(\position1/x_sum [11]), .B(n510), .Q(\position1/n1009 ) );
  NAND22 U2875 ( .A(\position1/N1188 ), .B(n638), .Q(\position1/n1011 ) );
  AOI221 U2876 ( .A(\position1/N496 ), .B(n740), .C(\position1/N915 ), .D(n640), .Q(\position1/n1010 ) );
  NAND41 U2877 ( .A(\position1/n1004 ), .B(\position1/n1005 ), .C(
        \position1/n1006 ), .D(\position1/n1007 ), .Q(\position1/n1623 ) );
  NAND22 U2878 ( .A(\position1/x_sum [12]), .B(n508), .Q(\position1/n1005 ) );
  NAND22 U2879 ( .A(\position1/N1189 ), .B(n635), .Q(\position1/n1007 ) );
  AOI221 U2880 ( .A(\position1/N497 ), .B(n740), .C(\position1/N916 ), .D(n639), .Q(\position1/n1006 ) );
  AOI221 U2881 ( .A(\position1/N342 ), .B(n644), .C(\position1/N619 ), .D(n645), .Q(\position1/n1004 ) );
  XOR21 U2882 ( .A(\position1/x_sum [12]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [12]), .Q(\position1/N619 )
         );
  XOR21 U2883 ( .A(\position1/N292 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [12]), .Q(
        \position1/N342 ) );
  NOR21 U2884 ( .A(n505), .B(\gensync1/N175 ), .Q(n2126) );
  XOR21 U2885 ( .A(\position1/y_sum [16]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [16]), .Q(\position1/N1218 )
         );
  XOR21 U2886 ( .A(\position1/x_sum [16]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [16]), .Q(\position1/N1193 )
         );
  XOR21 U2887 ( .A(\position1/y_sum [17]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [17]), .Q(\position1/N1219 )
         );
  XOR21 U2888 ( .A(\position1/x_sum [15]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [15]), .Q(\position1/N1192 )
         );
  AOI221 U2889 ( .A(\position1/N417 ), .B(n643), .C(\position1/N644 ), .D(n646), .Q(\position1/n904 ) );
  XOR21 U2890 ( .A(\position1/y_sum [12]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [12]), .Q(\position1/N644 )
         );
  XOR21 U2891 ( .A(\position1/N367 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [12]), .Q(
        \position1/N417 ) );
  AOI221 U2892 ( .A(\position1/N418 ), .B(n643), .C(\position1/N645 ), .D(n647), .Q(\position1/n900 ) );
  XOR21 U2893 ( .A(\position1/y_sum [13]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [13]), .Q(\position1/N645 )
         );
  XOR21 U2894 ( .A(\position1/N368 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [13]), .Q(
        \position1/N418 ) );
  AOI221 U2895 ( .A(\position1/N341 ), .B(n643), .C(\position1/N618 ), .D(n645), .Q(\position1/n1008 ) );
  XOR21 U2896 ( .A(\position1/x_sum [11]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [11]), .Q(\position1/N618 )
         );
  XOR21 U2897 ( .A(\position1/N291 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [11]), .Q(
        \position1/N341 ) );
  NAND41 U2898 ( .A(\position1/n912 ), .B(\position1/n913 ), .C(
        \position1/n914 ), .D(\position1/n915 ), .Q(\position1/n1600 ) );
  NAND22 U2899 ( .A(\position1/y_sum [10]), .B(n673), .Q(\position1/n913 ) );
  NAND22 U2900 ( .A(\position1/N1212 ), .B(n636), .Q(\position1/n915 ) );
  AOI221 U2901 ( .A(\position1/N415 ), .B(n643), .C(\position1/N642 ), .D(n645), .Q(\position1/n912 ) );
  NAND41 U2902 ( .A(\position1/n908 ), .B(\position1/n909 ), .C(
        \position1/n910 ), .D(\position1/n911 ), .Q(\position1/n1599 ) );
  NAND22 U2903 ( .A(\position1/y_sum [11]), .B(n509), .Q(\position1/n909 ) );
  NAND22 U2904 ( .A(\position1/N1213 ), .B(n637), .Q(\position1/n911 ) );
  AOI221 U2905 ( .A(\position1/N546 ), .B(n740), .C(\position1/N990 ), .D(n640), .Q(\position1/n910 ) );
  NAND41 U2906 ( .A(\position1/n1012 ), .B(\position1/n1013 ), .C(
        \position1/n1014 ), .D(\position1/n1015 ), .Q(\position1/n1625 ) );
  NAND22 U2907 ( .A(\position1/x_sum [10]), .B(n510), .Q(\position1/n1013 ) );
  NAND22 U2908 ( .A(\position1/N1187 ), .B(n638), .Q(\position1/n1015 ) );
  AOI221 U2909 ( .A(\position1/N495 ), .B(n740), .C(\position1/N914 ), .D(n641), .Q(\position1/n1014 ) );
  NAND41 U2910 ( .A(\position1/n916 ), .B(\position1/n917 ), .C(
        \position1/n918 ), .D(\position1/n919 ), .Q(\position1/n1601 ) );
  NAND22 U2911 ( .A(\position1/y_sum [9]), .B(n673), .Q(\position1/n917 ) );
  NAND22 U2912 ( .A(\position1/N1211 ), .B(n636), .Q(\position1/n919 ) );
  AOI221 U2913 ( .A(\position1/N544 ), .B(n740), .C(\position1/N988 ), .D(n640), .Q(\position1/n918 ) );
  NAND41 U2914 ( .A(\position1/n1020 ), .B(\position1/n1021 ), .C(
        \position1/n1022 ), .D(\position1/n1023 ), .Q(\position1/n1627 ) );
  NAND22 U2915 ( .A(\position1/x_sum [8]), .B(n510), .Q(\position1/n1021 ) );
  NAND22 U2916 ( .A(\position1/N1185 ), .B(n638), .Q(\position1/n1023 ) );
  AOI221 U2917 ( .A(\position1/N493 ), .B(n740), .C(\position1/N912 ), .D(
        \position1/n857 ), .Q(\position1/n1022 ) );
  NAND41 U2918 ( .A(\position1/n1016 ), .B(\position1/n1017 ), .C(
        \position1/n1018 ), .D(\position1/n1019 ), .Q(\position1/n1626 ) );
  NAND22 U2919 ( .A(\position1/x_sum [9]), .B(n510), .Q(\position1/n1017 ) );
  NAND22 U2920 ( .A(\position1/N1186 ), .B(n638), .Q(\position1/n1019 ) );
  AOI221 U2921 ( .A(\position1/N494 ), .B(n740), .C(\position1/N913 ), .D(
        \position1/n857 ), .Q(\position1/n1018 ) );
  AOI221 U2922 ( .A(\position1/N414 ), .B(n643), .C(\position1/N641 ), .D(n646), .Q(\position1/n916 ) );
  XOR21 U2923 ( .A(\position1/y_sum [9]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [9]), .Q(\position1/N641 )
         );
  AOI221 U2924 ( .A(\position1/N339 ), .B(n642), .C(\position1/N616 ), .D(n645), .Q(\position1/n1016 ) );
  XOR21 U2925 ( .A(\position1/x_sum [9]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [9]), .Q(\position1/N616 )
         );
  AOI221 U2926 ( .A(\position1/N340 ), .B(n644), .C(\position1/N617 ), .D(n645), .Q(\position1/n1012 ) );
  XOR21 U2927 ( .A(\position1/x_sum [10]), .B(
        \position1/dp_cluster_4/add_178_aco/carry [10]), .Q(\position1/N617 )
         );
  XOR21 U2928 ( .A(\position1/N290 ), .B(
        \position1/dp_cluster_7/add_0_root_add_170_3/carry [10]), .Q(
        \position1/N340 ) );
  XOR21 U2929 ( .A(\position1/y_sum [14]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [14]), .Q(\position1/N1216 )
         );
  XOR21 U2930 ( .A(\position1/x_sum [12]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [12]), .Q(\position1/N1189 )
         );
  XOR21 U2931 ( .A(\position1/x_sum [14]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [14]), .Q(\position1/N1191 )
         );
  XOR21 U2932 ( .A(\position1/y_sum [13]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [13]), .Q(\position1/N1215 )
         );
  XOR21 U2933 ( .A(\position1/y_sum [15]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [15]), .Q(\position1/N1217 )
         );
  XOR21 U2934 ( .A(\position1/x_sum [13]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [13]), .Q(\position1/N1190 )
         );
  AOI221 U2935 ( .A(\position1/N416 ), .B(n643), .C(\position1/N643 ), .D(n647), .Q(\position1/n908 ) );
  XOR21 U2936 ( .A(\position1/y_sum [11]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [11]), .Q(\position1/N643 )
         );
  XOR21 U2937 ( .A(\position1/N366 ), .B(
        \position1/dp_cluster_6/add_0_root_add_171_3/carry [11]), .Q(
        \position1/N416 ) );
  INV3 U2938 ( .A(\position1/n1153 ), .Q(n711) );
  AOI221 U2939 ( .A(\position1/N224 ), .B(n481), .C(\position1/count_img [19]), 
        .D(n483), .Q(\position1/n1153 ) );
  XOR21 U2940 ( .A(\position1/add_161/carry [19]), .B(
        \position1/count_img [19]), .Q(\position1/N224 ) );
  NAND41 U2941 ( .A(\position1/n924 ), .B(\position1/n925 ), .C(
        \position1/n926 ), .D(\position1/n927 ), .Q(\position1/n1603 ) );
  NAND22 U2942 ( .A(\position1/y_sum [7]), .B(n673), .Q(\position1/n925 ) );
  NAND22 U2943 ( .A(\position1/N1209 ), .B(n636), .Q(\position1/n927 ) );
  AOI221 U2944 ( .A(\position1/N542 ), .B(n740), .C(\position1/N986 ), .D(n640), .Q(\position1/n926 ) );
  NAND41 U2945 ( .A(\position1/n920 ), .B(\position1/n921 ), .C(
        \position1/n922 ), .D(\position1/n923 ), .Q(\position1/n1602 ) );
  NAND22 U2946 ( .A(\position1/y_sum [8]), .B(n673), .Q(\position1/n921 ) );
  NAND22 U2947 ( .A(\position1/N1210 ), .B(n636), .Q(\position1/n923 ) );
  AOI221 U2948 ( .A(\position1/N543 ), .B(n740), .C(\position1/N987 ), .D(n640), .Q(\position1/n922 ) );
  NAND41 U2949 ( .A(\position1/n1024 ), .B(\position1/n1025 ), .C(
        \position1/n1026 ), .D(\position1/n1027 ), .Q(\position1/n1628 ) );
  NAND22 U2950 ( .A(\position1/x_sum [7]), .B(n510), .Q(\position1/n1025 ) );
  NAND22 U2951 ( .A(\position1/N1184 ), .B(n638), .Q(\position1/n1027 ) );
  AOI221 U2952 ( .A(\position1/N492 ), .B(n740), .C(\position1/N911 ), .D(
        \position1/n857 ), .Q(\position1/n1026 ) );
  INV3 U2953 ( .A(\position1/n1157 ), .Q(n709) );
  AOI221 U2954 ( .A(\position1/N222 ), .B(\position1/n1154 ), .C(n482), .D(
        \position1/count_img [17]), .Q(\position1/n1157 ) );
  XOR21 U2955 ( .A(\position1/y_sum [12]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [12]), .Q(\position1/N1214 )
         );
  XOR21 U2956 ( .A(\position1/x_sum [10]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [10]), .Q(\position1/N1187 )
         );
  XOR21 U2957 ( .A(\position1/y_sum [11]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [11]), .Q(\position1/N1213 )
         );
  XOR21 U2958 ( .A(\position1/x_sum [11]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [11]), .Q(\position1/N1188 )
         );
  XOR21 U2959 ( .A(\position1/y_sum [10]), .B(
        \position1/dp_cluster_5/add_179_aco/carry [10]), .Q(\position1/N642 )
         );
  BUF2 U2960 ( .A(\position1/N560 ), .Q(n514) );
  BUF2 U2961 ( .A(\position1/N2460 ), .Q(n631) );
  BUF2 U2962 ( .A(\position1/N2459 ), .Q(n627) );
  INV3 U2963 ( .A(\position1/n1156 ), .Q(n710) );
  AOI221 U2964 ( .A(\position1/N223 ), .B(n480), .C(\position1/count_img [18]), 
        .D(n483), .Q(\position1/n1156 ) );
  NAND41 U2965 ( .A(\position1/n928 ), .B(\position1/n929 ), .C(
        \position1/n930 ), .D(\position1/n931 ), .Q(\position1/n1604 ) );
  NAND22 U2966 ( .A(\position1/y_sum [6]), .B(n673), .Q(\position1/n929 ) );
  NAND22 U2967 ( .A(\position1/N1208 ), .B(n636), .Q(\position1/n931 ) );
  AOI221 U2968 ( .A(\position1/N541 ), .B(n740), .C(\position1/N985 ), .D(n640), .Q(\position1/n930 ) );
  NAND41 U2969 ( .A(\position1/n1032 ), .B(\position1/n1033 ), .C(
        \position1/n1034 ), .D(\position1/n1035 ), .Q(\position1/n1630 ) );
  NAND22 U2970 ( .A(\position1/x_sum [5]), .B(n510), .Q(\position1/n1033 ) );
  NAND22 U2971 ( .A(\position1/N1182 ), .B(n638), .Q(\position1/n1035 ) );
  AOI221 U2972 ( .A(\position1/N490 ), .B(n740), .C(\position1/N909 ), .D(
        \position1/n857 ), .Q(\position1/n1034 ) );
  NAND41 U2973 ( .A(\position1/n1028 ), .B(\position1/n1029 ), .C(
        \position1/n1030 ), .D(\position1/n1031 ), .Q(\position1/n1629 ) );
  NAND22 U2974 ( .A(\position1/x_sum [6]), .B(n510), .Q(\position1/n1029 ) );
  NAND22 U2975 ( .A(\position1/N1183 ), .B(n638), .Q(\position1/n1031 ) );
  AOI221 U2976 ( .A(\position1/N491 ), .B(n740), .C(\position1/N910 ), .D(
        \position1/n857 ), .Q(\position1/n1030 ) );
  XOR21 U2977 ( .A(\position1/y_sum [10]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [10]), .Q(\position1/N1212 )
         );
  XOR21 U2978 ( .A(\position1/y_sum [9]), .B(
        \position1/dp_cluster_1/add_197_aco/carry [9]), .Q(\position1/N1211 )
         );
  XOR21 U2979 ( .A(\position1/x_sum [9]), .B(
        \position1/dp_cluster_0/add_196_aco/carry [9]), .Q(\position1/N1186 )
         );
  BUF2 U2980 ( .A(\position1/N2458 ), .Q(n623) );
  INV3 U2981 ( .A(\position1/n1158 ), .Q(n708) );
  AOI221 U2982 ( .A(\position1/N221 ), .B(n481), .C(n483), .D(
        \position1/count_img [16]), .Q(\position1/n1158 ) );
  NOR31 U2983 ( .A(n2125), .B(\position1/count_img [19]), .C(
        \position1/count_img [18]), .Q(\position1/N267 ) );
  AOI211 U2984 ( .A(n497), .B(\position1/n1390 ), .C(\position1/n1391 ), .Q(
        \position1/n1389 ) );
  NOR31 U2985 ( .A(n2124), .B(n2123), .C(n18), .Q(n2125) );
  NAND41 U2986 ( .A(\position1/N2402 ), .B(\position1/N2391 ), .C(
        \position1/N2413 ), .D(\position1/n1579 ), .Q(\position1/n1182 ) );
  NAND41 U2987 ( .A(\position1/n952 ), .B(\position1/n953 ), .C(
        \position1/n954 ), .D(\position1/n955 ), .Q(\position1/n1610 ) );
  NAND22 U2988 ( .A(\position1/N1938 ), .B(n673), .Q(\position1/n953 ) );
  AOI221 U2989 ( .A(\position1/N355 ), .B(n642), .C(\position1/N632 ), .D(n646), .Q(\position1/n952 ) );
  NAND22 U2990 ( .A(\position1/N1202 ), .B(n636), .Q(\position1/n955 ) );
  NAND41 U2991 ( .A(\position1/n1052 ), .B(\position1/n1053 ), .C(
        \position1/n1054 ), .D(\position1/n1055 ), .Q(\position1/n1635 ) );
  NAND22 U2992 ( .A(\position1/N1521 ), .B(n510), .Q(\position1/n1053 ) );
  AOI221 U2993 ( .A(\position1/N280 ), .B(\position1/n858 ), .C(
        \position1/N607 ), .D(n645), .Q(\position1/n1052 ) );
  NAND22 U2994 ( .A(\position1/N1177 ), .B(n638), .Q(\position1/n1055 ) );
  NAND41 U2995 ( .A(\position1/n948 ), .B(\position1/n949 ), .C(
        \position1/n950 ), .D(\position1/n951 ), .Q(\position1/n1609 ) );
  NAND22 U2996 ( .A(\position1/y_sum [1]), .B(n673), .Q(\position1/n949 ) );
  AOI221 U2997 ( .A(\position1/N406 ), .B(n643), .C(\position1/N633 ), .D(
        \position1/n859 ), .Q(\position1/n948 ) );
  NAND22 U2998 ( .A(\position1/N1203 ), .B(n636), .Q(\position1/n951 ) );
  NAND41 U2999 ( .A(\position1/n1048 ), .B(\position1/n1049 ), .C(
        \position1/n1050 ), .D(\position1/n1051 ), .Q(\position1/n1634 ) );
  NAND22 U3000 ( .A(\position1/x_sum [1]), .B(n510), .Q(\position1/n1049 ) );
  AOI221 U3001 ( .A(\position1/N331 ), .B(\position1/n858 ), .C(
        \position1/N608 ), .D(n645), .Q(\position1/n1048 ) );
  NAND22 U3002 ( .A(\position1/N1178 ), .B(n638), .Q(\position1/n1051 ) );
  NAND41 U3003 ( .A(\position1/n944 ), .B(\position1/n945 ), .C(
        \position1/n946 ), .D(\position1/n947 ), .Q(\position1/n1608 ) );
  NAND22 U3004 ( .A(\position1/y_sum [2]), .B(n673), .Q(\position1/n945 ) );
  AOI221 U3005 ( .A(\position1/N407 ), .B(n643), .C(\position1/N634 ), .D(
        \position1/n859 ), .Q(\position1/n944 ) );
  NAND22 U3006 ( .A(\position1/N1204 ), .B(n636), .Q(\position1/n947 ) );
  NAND41 U3007 ( .A(\position1/n940 ), .B(\position1/n941 ), .C(
        \position1/n942 ), .D(\position1/n943 ), .Q(\position1/n1607 ) );
  NAND22 U3008 ( .A(\position1/y_sum [3]), .B(n673), .Q(\position1/n941 ) );
  AOI221 U3009 ( .A(\position1/N408 ), .B(n643), .C(\position1/N635 ), .D(
        \position1/n859 ), .Q(\position1/n940 ) );
  NAND22 U3010 ( .A(\position1/N1205 ), .B(n636), .Q(\position1/n943 ) );
  NAND41 U3011 ( .A(\position1/n936 ), .B(\position1/n937 ), .C(
        \position1/n938 ), .D(\position1/n939 ), .Q(\position1/n1606 ) );
  NAND22 U3012 ( .A(\position1/y_sum [4]), .B(n673), .Q(\position1/n937 ) );
  AOI221 U3013 ( .A(\position1/N409 ), .B(n643), .C(\position1/N636 ), .D(
        \position1/n859 ), .Q(\position1/n936 ) );
  NAND22 U3014 ( .A(\position1/N1206 ), .B(n636), .Q(\position1/n939 ) );
  NAND41 U3015 ( .A(\position1/n932 ), .B(\position1/n933 ), .C(
        \position1/n934 ), .D(\position1/n935 ), .Q(\position1/n1605 ) );
  NAND22 U3016 ( .A(\position1/y_sum [5]), .B(n673), .Q(\position1/n933 ) );
  NAND22 U3017 ( .A(\position1/N1207 ), .B(n636), .Q(\position1/n935 ) );
  AOI221 U3018 ( .A(\position1/N410 ), .B(n643), .C(\position1/N637 ), .D(
        \position1/n859 ), .Q(\position1/n932 ) );
  NAND41 U3019 ( .A(\position1/n1044 ), .B(\position1/n1045 ), .C(
        \position1/n1046 ), .D(\position1/n1047 ), .Q(\position1/n1633 ) );
  NAND22 U3020 ( .A(\position1/x_sum [2]), .B(n510), .Q(\position1/n1045 ) );
  AOI221 U3021 ( .A(\position1/N332 ), .B(\position1/n858 ), .C(
        \position1/N609 ), .D(n645), .Q(\position1/n1044 ) );
  NAND22 U3022 ( .A(\position1/N1179 ), .B(n638), .Q(\position1/n1047 ) );
  NAND41 U3023 ( .A(\position1/n1040 ), .B(\position1/n1041 ), .C(
        \position1/n1042 ), .D(\position1/n1043 ), .Q(\position1/n1632 ) );
  NAND22 U3024 ( .A(\position1/x_sum [3]), .B(n673), .Q(\position1/n1041 ) );
  AOI221 U3025 ( .A(\position1/N333 ), .B(\position1/n858 ), .C(
        \position1/N610 ), .D(n645), .Q(\position1/n1040 ) );
  NAND22 U3026 ( .A(\position1/N1180 ), .B(n637), .Q(\position1/n1043 ) );
  NAND41 U3027 ( .A(\position1/n1036 ), .B(\position1/n1037 ), .C(
        \position1/n1038 ), .D(\position1/n1039 ), .Q(\position1/n1631 ) );
  NAND22 U3028 ( .A(\position1/x_sum [4]), .B(n673), .Q(\position1/n1037 ) );
  NAND22 U3029 ( .A(\position1/N1181 ), .B(n636), .Q(\position1/n1039 ) );
  AOI221 U3030 ( .A(\position1/N334 ), .B(\position1/n858 ), .C(
        \position1/N611 ), .D(n645), .Q(\position1/n1036 ) );
  INV3 U3031 ( .A(\position1/n1160 ), .Q(n706) );
  AOI221 U3032 ( .A(\position1/N219 ), .B(\position1/n1154 ), .C(
        \position1/count_img [14]), .D(n482), .Q(\position1/n1160 ) );
  AOI221 U3033 ( .A(n1389), .B(Y_barycentre_top[0]), .C(Y_barycentre_top[1]), 
        .D(\position1/N2383 ), .Q(n1391) );
  AOI211 U3034 ( .A(\position1/N2405 ), .B(n23), .C(\gensync1/n99 ), .Q(n1389)
         );
  XNR21 U3035 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [2]), 
        .B(cam_y[0]), .Q(\position1/N2405 ) );
  NOR21 U3036 ( .A(X_barycentre_top[6]), .B(n846), .Q(n1444) );
  INV3 U3037 ( .A(\position1/N2378 ), .Q(n846) );
  INV3 U3038 ( .A(\position1/n1178 ), .Q(n715) );
  AOI211 U3039 ( .A(reset_top), .B(\position1/gi [7]), .C(\position1/n1179 ), 
        .Q(\position1/n1178 ) );
  INV3 U3040 ( .A(\position1/n1180 ), .Q(n714) );
  AOI211 U3041 ( .A(reset_top), .B(\position1/gi [3]), .C(\position1/n1179 ), 
        .Q(\position1/n1180 ) );
  INV3 U3042 ( .A(\position1/n1181 ), .Q(n713) );
  AOI211 U3043 ( .A(reset_top), .B(\position1/gi [1]), .C(\position1/n1179 ), 
        .Q(\position1/n1181 ) );
  AOI2111 U3044 ( .A(\position1/n1580 ), .B(\position1/n1581 ), .C(n843), .D(
        \position1/n1582 ), .Q(\position1/n1579 ) );
  NOR40 U3045 ( .A(Y_barycentre_top[3]), .B(Y_barycentre_top[2]), .C(
        Y_barycentre_top[1]), .D(Y_barycentre_top[0]), .Q(\position1/n1580 )
         );
  NOR40 U3046 ( .A(Y_barycentre_top[6]), .B(n878), .C(Y_barycentre_top[5]), 
        .D(Y_barycentre_top[4]), .Q(\position1/n1581 ) );
  NOR40 U3047 ( .A(n879), .B(n880), .C(X_barycentre_top[5]), .D(
        X_barycentre_top[4]), .Q(\position1/n1582 ) );
  NOR21 U3048 ( .A(\position1/n1177 ), .B(\position1/n368 ), .Q(
        \position1/N99 ) );
  NOR21 U3049 ( .A(\position1/n1177 ), .B(\position1/n369 ), .Q(
        \position1/N98 ) );
  NOR21 U3050 ( .A(\position1/n1177 ), .B(\position1/n370 ), .Q(
        \position1/N97 ) );
  NOR21 U3051 ( .A(\position1/n1177 ), .B(\position1/n346 ), .Q(
        \position1/N88 ) );
  NOR21 U3052 ( .A(\position1/n1177 ), .B(\position1/n347 ), .Q(
        \position1/N87 ) );
  NOR21 U3053 ( .A(\position1/n1177 ), .B(\position1/n348 ), .Q(
        \position1/N86 ) );
  NOR21 U3054 ( .A(\position1/n1177 ), .B(\position1/n349 ), .Q(
        \position1/N85 ) );
  NOR21 U3055 ( .A(\position1/n1177 ), .B(\position1/n350 ), .Q(
        \position1/N84 ) );
  NOR21 U3056 ( .A(\position1/n1177 ), .B(\position1/n351 ), .Q(
        \position1/N83 ) );
  NOR21 U3057 ( .A(\position1/n1177 ), .B(\position1/n352 ), .Q(
        \position1/N82 ) );
  NOR21 U3058 ( .A(\position1/n1177 ), .B(\position1/n353 ), .Q(
        \position1/N81 ) );
  NOR21 U3059 ( .A(\position1/n1177 ), .B(\position1/n363 ), .Q(
        \position1/N104 ) );
  NOR21 U3060 ( .A(\position1/n1177 ), .B(\position1/n364 ), .Q(
        \position1/N103 ) );
  NOR21 U3061 ( .A(\position1/n1177 ), .B(\position1/n365 ), .Q(
        \position1/N102 ) );
  NOR21 U3062 ( .A(\position1/n1177 ), .B(\position1/n366 ), .Q(
        \position1/N101 ) );
  NOR21 U3063 ( .A(\position1/n1177 ), .B(\position1/n367 ), .Q(
        \position1/N100 ) );
  AOI221 U3064 ( .A(\position1/N2395 ), .B(n16), .C(n1406), .D(n1405), .Q(
        n1407) );
  INV3 U3065 ( .A(\position1/N2396 ), .Q(n841) );
  AOI221 U3066 ( .A(Y_barycentre_top[2]), .B(n806), .C(n1421), .D(n1420), .Q(
        n1422) );
  NAND22 U3067 ( .A(\position1/N2384 ), .B(n21), .Q(n1420) );
  INV3 U3068 ( .A(\position1/N2384 ), .Q(n806) );
  AOI221 U3069 ( .A(n1419), .B(\gensync1/n99 ), .C(\position1/N2383 ), .D(n23), 
        .Q(n1421) );
  AOI221 U3070 ( .A(n1434), .B(n211), .C(\position1/N2373 ), .D(n17), .Q(n1436) );
  AOI211 U3071 ( .A(X_barycentre_top[1]), .B(\position1/N2394 ), .C(
        X_barycentre_top[0]), .Q(n1434) );
  XOR21 U3072 ( .A(n501), .B(cam_x[0]), .Q(\position1/N2373 ) );
  AOI221 U3073 ( .A(X_barycentre_top[2]), .B(n850), .C(n1436), .D(n1435), .Q(
        n1437) );
  NAND22 U3074 ( .A(\position1/N2374 ), .B(n16), .Q(n1435) );
  INV3 U3075 ( .A(\position1/N2374 ), .Q(n850) );
  INV3 U3076 ( .A(\position1/N2385 ), .Q(n802) );
  XNR21 U3077 ( .A(\position1/dp_cluster_6/add_1_root_add_171_3/carry [4]), 
        .B(\position1/sub_250_3/carry[3] ), .Q(\position1/N2385 ) );
  NOR21 U3078 ( .A(Y_barycentre_top[7]), .B(n785), .Q(n1401) );
  NOR21 U3079 ( .A(\position1/N2410 ), .B(n31), .Q(n1399) );
  AOI221 U3080 ( .A(n1404), .B(X_barycentre_top[0]), .C(X_barycentre_top[1]), 
        .D(\position1/N2373 ), .Q(n1406) );
  AOI211 U3081 ( .A(\position1/N2394 ), .B(n17), .C(n211), .Q(n1404) );
  XNR21 U3082 ( .A(n501), .B(cam_x[0]), .Q(\position1/N2394 ) );
  NOR21 U3083 ( .A(X_barycentre_top[5]), .B(n839), .Q(n1412) );
  NOR21 U3084 ( .A(\position1/N2397 ), .B(n20), .Q(n1410) );
  NOR21 U3085 ( .A(Y_barycentre_top[5]), .B(n793), .Q(n1397) );
  NOR21 U3086 ( .A(\position1/N2408 ), .B(n26), .Q(n1395) );
  NOR21 U3087 ( .A(X_barycentre_top[4]), .B(n848), .Q(n1440) );
  INV3 U3088 ( .A(\position1/N2375 ), .Q(n849) );
  NOR21 U3089 ( .A(Y_barycentre_top[4]), .B(n798), .Q(n1425) );
  INV3 U3090 ( .A(\position1/N2386 ), .Q(n798) );
  NOR21 U3091 ( .A(X_barycentre_top[7]), .B(n837), .Q(n1416) );
  NOR21 U3092 ( .A(\position1/N2399 ), .B(n25), .Q(n1414) );
  BUF2 U3093 ( .A(\position1/N2456 ), .Q(n620) );
  INV3 U3094 ( .A(\position1/N2387 ), .Q(n794) );
  NOR21 U3095 ( .A(\position1/N2387 ), .B(n28), .Q(n1427) );
  INV3 U3096 ( .A(\position1/N2389 ), .Q(n786) );
  NOR21 U3097 ( .A(\position1/N2389 ), .B(n32), .Q(n1431) );
  NAND22 U3098 ( .A(X_barycentre_top[2]), .B(n842), .Q(n1405) );
  INV3 U3099 ( .A(\position1/N2395 ), .Q(n842) );
  NAND22 U3100 ( .A(Y_barycentre_top[2]), .B(n805), .Q(n1390) );
  INV3 U3101 ( .A(\position1/N2406 ), .Q(n805) );
  NOR21 U3102 ( .A(Y_barycentre_top[8]), .B(n780), .Q(n1433) );
  INV3 U3103 ( .A(\position1/N2390 ), .Q(n780) );
  NOR21 U3104 ( .A(Y_barycentre_top[6]), .B(n790), .Q(n1429) );
  INV3 U3105 ( .A(\position1/N2388 ), .Q(n790) );
  AOI221 U3106 ( .A(\position1/N2406 ), .B(n21), .C(n1391), .D(n1390), .Q(
        n1392) );
  INV3 U3107 ( .A(\position1/N2407 ), .Q(n801) );
  INV3 U3108 ( .A(\position1/N2381 ), .Q(n843) );
  NOR21 U3109 ( .A(X_barycentre_top[8]), .B(n844), .Q(n1448) );
  AOI211 U3110 ( .A(Y_barycentre_top[1]), .B(\position1/N2405 ), .C(
        Y_barycentre_top[0]), .Q(n1419) );
  INV3 U3111 ( .A(\position1/n1159 ), .Q(n707) );
  AOI221 U3112 ( .A(\position1/N220 ), .B(n480), .C(n483), .D(
        \position1/count_img [15]), .Q(\position1/n1159 ) );
  BUF2 U3113 ( .A(\position1/N2460 ), .Q(n630) );
  BUF2 U3114 ( .A(\position1/N2455 ), .Q(n469) );
  BUF2 U3115 ( .A(\position1/N560 ), .Q(n515) );
  BUF2 U3116 ( .A(\position1/N2454 ), .Q(n615) );
  INV3 U3117 ( .A(\position1/n1162 ), .Q(n704) );
  AOI221 U3118 ( .A(\position1/N217 ), .B(n480), .C(\position1/count_img [12]), 
        .D(n483), .Q(\position1/n1162 ) );
  INV3 U3119 ( .A(\position1/n1161 ), .Q(n705) );
  AOI221 U3120 ( .A(\position1/N218 ), .B(n481), .C(n483), .D(
        \position1/count_img [13]), .Q(\position1/n1161 ) );
  INV3 U3121 ( .A(\position1/n1163 ), .Q(n703) );
  AOI221 U3122 ( .A(\position1/N216 ), .B(\position1/n1154 ), .C(n482), .D(
        \position1/count_img [11]), .Q(\position1/n1163 ) );
  BUF2 U3123 ( .A(\position1/N2458 ), .Q(n621) );
  BUF2 U3124 ( .A(\position1/N2459 ), .Q(n625) );
  AOI211 U3125 ( .A(\image_process1/n91 ), .B(\image_process1/gi [7]), .C(
        \image_process1/n89 ), .Q(\image_process1/n86 ) );
  AOI211 U3126 ( .A(\image_process1/n91 ), .B(\image_process1/gi [3]), .C(
        \image_process1/n89 ), .Q(\image_process1/n106 ) );
  AOI211 U3127 ( .A(\image_process1/n91 ), .B(\image_process1/gi [1]), .C(
        \image_process1/n89 ), .Q(\image_process1/n114 ) );
  INV3 U3128 ( .A(\image_process1/n88 ), .Q(n772) );
  AOI211 U3129 ( .A(\image_process1/n58 ), .B(\image_process1/gi [7]), .C(
        \image_process1/n89 ), .Q(\image_process1/n88 ) );
  INV3 U3130 ( .A(\image_process1/n108 ), .Q(n768) );
  AOI211 U3131 ( .A(\image_process1/n58 ), .B(\image_process1/gi [3]), .C(
        \image_process1/n89 ), .Q(\image_process1/n108 ) );
  INV3 U3132 ( .A(\image_process1/n116 ), .Q(n766) );
  AOI211 U3133 ( .A(\image_process1/n58 ), .B(\image_process1/gi [1]), .C(
        \image_process1/n89 ), .Q(\image_process1/n116 ) );
  AOI211 U3134 ( .A(\position1/count_img [13]), .B(n1353), .C(
        \position1/count_img [14]), .Q(n2123) );
  INV3 U3135 ( .A(n2122), .Q(n1353) );
  AOI311 U3136 ( .A(\position1/count_img [10]), .B(n1354), .C(
        \position1/count_img [11]), .D(\position1/count_img [12]), .Q(n2122)
         );
  INV3 U3137 ( .A(n2121), .Q(n1354) );
  AOI211 U3138 ( .A(\position1/count_img [8]), .B(n2120), .C(
        \position1/count_img [9]), .Q(n2121) );
  NOR21 U3139 ( .A(\position1/count_img [7]), .B(\position1/count_img [6]), 
        .Q(n2117) );
  NAND31 U3140 ( .A(\position1/count_img [1]), .B(\position1/count_img [0]), 
        .C(\position1/count_img [2]), .Q(n2119) );
  NAND31 U3141 ( .A(\position1/count_img [4]), .B(\position1/count_img [3]), 
        .C(\position1/count_img [5]), .Q(n2118) );
  XNR21 U3142 ( .A(\gensync1/add_45/carry [9]), .B(\gensync1/comptY[9] ), .Q(
        n112) );
  BUF2 U3143 ( .A(\position1/N2455 ), .Q(n470) );
  BUF2 U3144 ( .A(\position1/N2456 ), .Q(n618) );
  BUF2 U3145 ( .A(\position1/N2452 ), .Q(n608) );
  NAND22 U3146 ( .A(\image_process1/n86 ), .B(\image_process1/n87 ), .Q(
        \image_process1/N31 ) );
  NAND22 U3147 ( .A(\image_process1/bi [7]), .B(n488), .Q(\image_process1/n87 ) );
  NAND22 U3148 ( .A(\image_process1/n106 ), .B(\image_process1/n107 ), .Q(
        \image_process1/N19 ) );
  NAND22 U3149 ( .A(\image_process1/bi [3]), .B(n488), .Q(
        \image_process1/n107 ) );
  NAND22 U3150 ( .A(\image_process1/n114 ), .B(\image_process1/n115 ), .Q(
        \image_process1/N13 ) );
  NAND22 U3151 ( .A(\image_process1/bi [1]), .B(n488), .Q(
        \image_process1/n115 ) );
  NAND22 U3152 ( .A(\image_process1/n86 ), .B(\image_process1/n90 ), .Q(
        \image_process1/N29 ) );
  NAND22 U3153 ( .A(\image_process1/ri [7]), .B(n488), .Q(\image_process1/n90 ) );
  NAND22 U3154 ( .A(\image_process1/n106 ), .B(\image_process1/n109 ), .Q(
        \image_process1/N17 ) );
  NAND22 U3155 ( .A(\image_process1/ri [3]), .B(n488), .Q(
        \image_process1/n109 ) );
  NAND22 U3156 ( .A(\image_process1/n114 ), .B(\image_process1/n118 ), .Q(
        \image_process1/N11 ) );
  NAND22 U3157 ( .A(\image_process1/ri [1]), .B(n488), .Q(
        \image_process1/n118 ) );
  INV3 U3158 ( .A(\position1/n1165 ), .Q(n701) );
  AOI221 U3159 ( .A(\position1/N214 ), .B(n480), .C(\position1/count_img [9]), 
        .D(n483), .Q(\position1/n1165 ) );
  INV3 U3160 ( .A(\position1/n1164 ), .Q(n702) );
  AOI221 U3161 ( .A(\position1/N215 ), .B(n481), .C(n483), .D(
        \position1/count_img [10]), .Q(\position1/n1164 ) );
  NOR31 U3162 ( .A(\image_process1/n27 ), .B(SW1_top), .C(\gensync1/n103 ), 
        .Q(\image_process1/n91 ) );
  AOI221 U3163 ( .A(\image_process1/n56 ), .B(\image_process1/n57 ), .C(
        \image_process1/gi [0]), .D(\image_process1/n91 ), .Q(
        \image_process1/n59 ) );
  AOI211 U3164 ( .A(\image_process1/n91 ), .B(\image_process1/gi [6]), .C(
        \image_process1/n95 ), .Q(\image_process1/n92 ) );
  AOI211 U3165 ( .A(\image_process1/n91 ), .B(\image_process1/gi [5]), .C(n776), .Q(\image_process1/n98 ) );
  AOI211 U3166 ( .A(\image_process1/n91 ), .B(\image_process1/gi [4]), .C(n776), .Q(\image_process1/n102 ) );
  AOI221 U3167 ( .A(\image_process1/n57 ), .B(\image_process1/n112 ), .C(
        \image_process1/n91 ), .D(\image_process1/gi [2]), .Q(
        \image_process1/n110 ) );
  NOR21 U3168 ( .A(\gensync1/n103 ), .B(\image_process1/state ), .Q(
        \image_process1/n61 ) );
  INV3 U3169 ( .A(\image_process1/n111 ), .Q(n767) );
  AOI221 U3170 ( .A(\image_process1/n57 ), .B(\image_process1/n112 ), .C(
        \image_process1/n58 ), .D(\image_process1/gi [2]), .Q(
        \image_process1/n111 ) );
  XNR21 U3171 ( .A(\gensync1/add_39/carry [9]), .B(\gensync1/N174 ), .Q(n113)
         );
  BUF2 U3172 ( .A(\position1/N2452 ), .Q(n607) );
  XOR21 U3173 ( .A(\position1/N1938 ), .B(n809), .Q(\position1/N632 ) );
  XOR21 U3174 ( .A(\position1/N1521 ), .B(n852), .Q(\position1/N607 ) );
  BUF2 U3175 ( .A(\position1/N2454 ), .Q(n613) );
  BUF2 U3176 ( .A(\position1/N2451 ), .Q(n473) );
  BUF2 U3177 ( .A(\position1/N2450 ), .Q(n605) );
  NAND22 U3178 ( .A(\image_process1/n92 ), .B(\image_process1/n93 ), .Q(
        \image_process1/N28 ) );
  NAND22 U3179 ( .A(\image_process1/bi [6]), .B(n488), .Q(\image_process1/n93 ) );
  NAND22 U3180 ( .A(\image_process1/n98 ), .B(\image_process1/n99 ), .Q(
        \image_process1/N25 ) );
  NAND22 U3181 ( .A(\image_process1/bi [5]), .B(n488), .Q(\image_process1/n99 ) );
  NAND22 U3182 ( .A(\image_process1/n102 ), .B(\image_process1/n103 ), .Q(
        \image_process1/N22 ) );
  NAND22 U3183 ( .A(\image_process1/bi [4]), .B(n488), .Q(
        \image_process1/n103 ) );
  NAND22 U3184 ( .A(\image_process1/n92 ), .B(\image_process1/n96 ), .Q(
        \image_process1/N26 ) );
  NAND22 U3185 ( .A(\image_process1/ri [6]), .B(n488), .Q(\image_process1/n96 ) );
  NAND22 U3186 ( .A(\image_process1/n98 ), .B(\image_process1/n101 ), .Q(
        \image_process1/N23 ) );
  NAND22 U3187 ( .A(\image_process1/ri [5]), .B(n488), .Q(
        \image_process1/n101 ) );
  NAND22 U3188 ( .A(\image_process1/n102 ), .B(\image_process1/n105 ), .Q(
        \image_process1/N20 ) );
  NAND22 U3189 ( .A(\image_process1/ri [4]), .B(n488), .Q(
        \image_process1/n105 ) );
  NAND22 U3190 ( .A(\image_process1/n59 ), .B(\image_process1/n119 ), .Q(
        \image_process1/N10 ) );
  NAND22 U3191 ( .A(\image_process1/bi [0]), .B(n488), .Q(
        \image_process1/n119 ) );
  NAND22 U3192 ( .A(\image_process1/n59 ), .B(\image_process1/n60 ), .Q(
        \image_process1/N8 ) );
  NAND22 U3193 ( .A(\image_process1/ri [0]), .B(n488), .Q(\image_process1/n60 ) );
  INV3 U3194 ( .A(\image_process1/n55 ), .Q(n773) );
  AOI221 U3195 ( .A(\image_process1/n56 ), .B(\image_process1/n57 ), .C(
        \image_process1/n58 ), .D(\image_process1/gi [0]), .Q(
        \image_process1/n55 ) );
  INV3 U3196 ( .A(\image_process1/n100 ), .Q(n770) );
  AOI211 U3197 ( .A(\image_process1/n58 ), .B(\image_process1/gi [5]), .C(n776), .Q(\image_process1/n100 ) );
  INV3 U3198 ( .A(\image_process1/n104 ), .Q(n769) );
  AOI211 U3199 ( .A(\image_process1/n58 ), .B(\image_process1/gi [4]), .C(n776), .Q(\image_process1/n104 ) );
  INV3 U3200 ( .A(\image_process1/n94 ), .Q(n771) );
  AOI211 U3201 ( .A(\image_process1/n58 ), .B(\image_process1/gi [6]), .C(
        \image_process1/n95 ), .Q(\image_process1/n94 ) );
  INV3 U3202 ( .A(\position1/n1174 ), .Q(n692) );
  AOI221 U3203 ( .A(\position1/n802 ), .B(n480), .C(n483), .D(
        \position1/count_img [0]), .Q(\position1/n1174 ) );
  INV3 U3204 ( .A(\position1/n1173 ), .Q(n693) );
  AOI221 U3205 ( .A(\position1/N206 ), .B(n481), .C(n483), .D(
        \position1/count_img [1]), .Q(\position1/n1173 ) );
  INV3 U3206 ( .A(\position1/n1171 ), .Q(n695) );
  AOI221 U3207 ( .A(\position1/N208 ), .B(n480), .C(n482), .D(
        \position1/count_img [3]), .Q(\position1/n1171 ) );
  INV3 U3208 ( .A(\position1/n1170 ), .Q(n696) );
  AOI221 U3209 ( .A(\position1/N209 ), .B(n481), .C(n482), .D(
        \position1/count_img [4]), .Q(\position1/n1170 ) );
  INV3 U3210 ( .A(\position1/n1168 ), .Q(n698) );
  AOI221 U3211 ( .A(\position1/N211 ), .B(n480), .C(\position1/count_img [6]), 
        .D(n483), .Q(\position1/n1168 ) );
  INV3 U3212 ( .A(\position1/n1167 ), .Q(n699) );
  AOI221 U3213 ( .A(\position1/N212 ), .B(n481), .C(\position1/count_img [7]), 
        .D(n483), .Q(\position1/n1167 ) );
  INV3 U3214 ( .A(\position1/n1172 ), .Q(n694) );
  AOI221 U3215 ( .A(\position1/N207 ), .B(\position1/n1154 ), .C(n483), .D(
        \position1/count_img [2]), .Q(\position1/n1172 ) );
  INV3 U3216 ( .A(\position1/n1169 ), .Q(n697) );
  AOI221 U3217 ( .A(\position1/N210 ), .B(\position1/n1154 ), .C(n483), .D(
        \position1/count_img [5]), .Q(\position1/n1169 ) );
  INV3 U3218 ( .A(\position1/n1166 ), .Q(n700) );
  AOI221 U3219 ( .A(\position1/N213 ), .B(\position1/n1154 ), .C(n483), .D(
        \position1/count_img [8]), .Q(\position1/n1166 ) );
  NOR40 U3220 ( .A(\position1/n1401 ), .B(\position1/n1402 ), .C(n1352), .D(
        n1350), .Q(\position1/n1144 ) );
  INV3 U3221 ( .A(\position1/n1403 ), .Q(n1350) );
  INV3 U3222 ( .A(\position1/n1405 ), .Q(n1352) );
  NAND41 U3223 ( .A(n1351), .B(\position1/count_img [16]), .C(
        \position1/count_img [13]), .D(\position1/count_img [15]), .Q(
        \position1/n1402 ) );
  NAND41 U3224 ( .A(n1356), .B(\position1/count_img [4]), .C(
        \position1/count_img [2]), .D(\position1/count_img [3]), .Q(
        \position1/n1401 ) );
  INV3 U3225 ( .A(\position1/n1408 ), .Q(n1356) );
  NAND22 U3226 ( .A(\position1/count_img [8]), .B(\position1/count_img [5]), 
        .Q(\position1/n1408 ) );
  NOR40 U3227 ( .A(\position1/n1406 ), .B(\position1/n802 ), .C(
        \position1/count_img [14]), .D(\position1/count_img [12]), .Q(
        \position1/n1405 ) );
  NAND22 U3228 ( .A(\position1/count_img [11]), .B(\position1/count_img [10]), 
        .Q(\position1/n1406 ) );
  XOR21 U3229 ( .A(\position1/N1938 ), .B(n810), .Q(\position1/N1202 ) );
  XOR21 U3230 ( .A(\position1/N1521 ), .B(n853), .Q(\position1/N1177 ) );
  BUF2 U3231 ( .A(\position1/N2451 ), .Q(n472) );
  BUF2 U3232 ( .A(\position1/N2450 ), .Q(n604) );
  BUF2 U3233 ( .A(\position1/N2448 ), .Q(n601) );
  NOR40 U3234 ( .A(\position1/count_img [6]), .B(n1355), .C(
        \position1/count_img [19]), .D(\position1/count_img [18]), .Q(
        \position1/n1403 ) );
  INV3 U3235 ( .A(\position1/n1404 ), .Q(n1355) );
  NOR21 U3236 ( .A(\position1/count_img [7]), .B(\position1/count_img [9]), 
        .Q(\position1/n1404 ) );
  NAND22 U3237 ( .A(\position1/count_img [17]), .B(\position1/count_img [16]), 
        .Q(n2124) );
  INV3 U3238 ( .A(\position1/n1407 ), .Q(n1351) );
  NAND22 U3239 ( .A(\position1/count_img [1]), .B(\position1/count_img [17]), 
        .Q(\position1/n1407 ) );
  AOI2111 U3240 ( .A(\image_process1/gi [5]), .B(n877), .C(
        \image_process1/gi [7]), .D(\image_process1/gi [6]), .Q(
        \image_process1/N62 ) );
  INV3 U3241 ( .A(n1386), .Q(n877) );
  AOI2111 U3242 ( .A(\image_process1/gi [2]), .B(\image_process1/gi [1]), .C(
        \image_process1/gi [4]), .D(\image_process1/gi [3]), .Q(n1386) );
  NOR40 U3243 ( .A(\position1/gi [2]), .B(\position1/gi [4]), .C(
        \position1/gi [5]), .D(\position1/gi [6]), .Q(\position1/n1148 ) );
  NAND31 U3244 ( .A(\position1/n1147 ), .B(\position1/n362 ), .C(
        \position1/n1148 ), .Q(\position1/n1058 ) );
  AOI211 U3245 ( .A(\image_process1/gi [6]), .B(n1385), .C(
        \image_process1/gi [7]), .Q(\image_process1/N64 ) );
  NOR40 U3246 ( .A(\image_process1/gi [3]), .B(\image_process1/gi [2]), .C(
        \image_process1/gi [1]), .D(\image_process1/gi [0]), .Q(n1384) );
  NAND31 U3247 ( .A(\position1/n1147 ), .B(\position1/gi [0]), .C(
        \position1/n1148 ), .Q(\position1/n1065 ) );
  NOR40 U3248 ( .A(\position1/n357 ), .B(\position1/n360 ), .C(
        \position1/n362 ), .D(\position1/gi [6]), .Q(\position1/n1150 ) );
  NAND31 U3249 ( .A(\position1/n1150 ), .B(\position1/n358 ), .C(
        \position1/n1147 ), .Q(\position1/n1146 ) );
  NAND31 U3250 ( .A(\position1/n1147 ), .B(\position1/n1150 ), .C(
        \position1/gi [4]), .Q(\position1/n1149 ) );
  NOR21 U3251 ( .A(\position1/n344 ), .B(\position1/state [0]), .Q(
        \position1/n1176 ) );
  BUF2 U3252 ( .A(\position1/N2448 ), .Q(n600) );
  NAND22 U3253 ( .A(\position1/state [1]), .B(\position1/state [0]), .Q(
        \position1/n1152 ) );
  INV3 U3254 ( .A(reset_top), .Q(n654) );
  NAND22 U3255 ( .A(n1387), .B(n5), .Q(n1388) );
  OAI311 U3256 ( .A(\image_process1/gi [0]), .B(\image_process1/gi [2]), .C(
        \image_process1/gi [1]), .D(\image_process1/gi [3]), .Q(n1387) );
  INV3 U3257 ( .A(\position1/n1584 ), .Q(n879) );
  NOR40 U3258 ( .A(X_barycentre_top[0]), .B(X_barycentre_top[1]), .C(
        X_barycentre_top[2]), .D(X_barycentre_top[3]), .Q(\position1/n1584 )
         );
  INV3 U3259 ( .A(\position1/n1583 ), .Q(n880) );
  NOR31 U3260 ( .A(X_barycentre_top[7]), .B(X_barycentre_top[8]), .C(
        X_barycentre_top[6]), .Q(\position1/n1583 ) );
  NOR31 U3261 ( .A(\gensync1/N167 ), .B(\gensync1/N165 ), .C(\gensync1/N166 ), 
        .Q(n1372) );
  OAI311 U3262 ( .A(\gensync1/N173 ), .B(\gensync1/N171 ), .C(\gensync1/N172 ), 
        .D(\gensync1/N170 ), .Q(n1373) );
  NOR31 U3263 ( .A(\gensync1/N181 ), .B(\gensync1/N74 ), .C(\gensync1/N182 ), 
        .Q(\gensync1/n90 ) );
  NAND22 U3264 ( .A(\image_process1/state ), .B(SW1_top), .Q(
        \image_process1/n117 ) );
  NOR21 U3265 ( .A(n506), .B(\gensync1/N173 ), .Q(\gensync1/N56 ) );
  BUF2 U3266 ( .A(\position1/N2445 ), .Q(n592) );
  BUF2 U3267 ( .A(\position1/N2446 ), .Q(n596) );
  NOR41 U3268 ( .A(\gensync1/n87 ), .B(n873), .C(\gensync1/N175 ), .D(
        \gensync1/N174 ), .Q(\gensync1/n107 ) );
  INV3 U3269 ( .A(\gensync1/n88 ), .Q(n873) );
  NAND22 U3270 ( .A(\gensync1/n89 ), .B(\gensync1/n90 ), .Q(\gensync1/n87 ) );
  NOR31 U3271 ( .A(\gensync1/N176 ), .B(\gensync1/N178 ), .C(\gensync1/N177 ), 
        .Q(\gensync1/n88 ) );
  BUF2 U3272 ( .A(\position1/N2446 ), .Q(n597) );
  NAND22 U3273 ( .A(reset_top), .B(\gensync1/N43 ), .Q(\gensync1/n101 ) );
  NAND22 U3274 ( .A(\gensync1/comptY[9] ), .B(n1375), .Q(\gensync1/N43 ) );
  NAND31 U3275 ( .A(n1374), .B(n1373), .C(n1372), .Q(n1375) );
  NOR21 U3276 ( .A(\gensync1/N168 ), .B(\gensync1/N169 ), .Q(n1374) );
  INV3 U3277 ( .A(reset_top), .Q(n650) );
  BUF2 U3278 ( .A(\position1/N2445 ), .Q(n594) );
  INV3 U3279 ( .A(\position1/n1585 ), .Q(n878) );
  NOR21 U3280 ( .A(Y_barycentre_top[7]), .B(Y_barycentre_top[8]), .Q(
        \position1/n1585 ) );
  INV3 U3281 ( .A(\position1/N2353 ), .Q(n1358) );
  INV3 U3282 ( .A(\position1/n843 ), .Q(n682) );
  AOI221 U3283 ( .A(n484), .B(X_barycentre_top[8]), .C(n634), .D(
        \position1/quot_x [8]), .Q(\position1/n843 ) );
  INV3 U3284 ( .A(\position1/n845 ), .Q(n680) );
  AOI221 U3285 ( .A(n484), .B(X_barycentre_top[6]), .C(n634), .D(
        \position1/quot_x [6]), .Q(\position1/n845 ) );
  INV3 U3286 ( .A(\position1/n844 ), .Q(n681) );
  AOI221 U3287 ( .A(n484), .B(X_barycentre_top[7]), .C(n634), .D(
        \position1/quot_x [7]), .Q(\position1/n844 ) );
  INV3 U3288 ( .A(\position1/n848 ), .Q(n677) );
  AOI221 U3289 ( .A(n484), .B(X_barycentre_top[3]), .C(n634), .D(
        \position1/quot_x [3]), .Q(\position1/n848 ) );
  INV3 U3290 ( .A(\position1/n849 ), .Q(n676) );
  AOI221 U3291 ( .A(n484), .B(X_barycentre_top[2]), .C(n634), .D(
        \position1/quot_x [2]), .Q(\position1/n849 ) );
  INV3 U3292 ( .A(\position1/n841 ), .Q(n684) );
  AOI221 U3293 ( .A(n484), .B(Y_barycentre_top[1]), .C(n634), .D(
        \position1/quot_y [1]), .Q(\position1/n841 ) );
  INV3 U3294 ( .A(\position1/n850 ), .Q(n675) );
  AOI221 U3295 ( .A(n484), .B(X_barycentre_top[1]), .C(n634), .D(
        \position1/quot_x [1]), .Q(\position1/n850 ) );
  INV3 U3296 ( .A(\position1/n842 ), .Q(n683) );
  AOI221 U3297 ( .A(n484), .B(Y_barycentre_top[0]), .C(n634), .D(
        \position1/quot_y [0]), .Q(\position1/n842 ) );
  INV3 U3298 ( .A(\position1/n851 ), .Q(n674) );
  AOI221 U3299 ( .A(n484), .B(X_barycentre_top[0]), .C(n633), .D(
        \position1/quot_x [0]), .Q(\position1/n851 ) );
  AOI211 U3300 ( .A(n1357), .B(\position1/n1383 ), .C(n652), .Q(
        \position1/N194 ) );
  NAND22 U3301 ( .A(\position1/n344 ), .B(\position1/state [0]), .Q(
        \position1/n1383 ) );
  INV3 U3302 ( .A(\position1/n1176 ), .Q(n1357) );
  OAI2111 U3303 ( .A(\gensync1/N178 ), .B(n874), .C(\gensync1/N175 ), .D(
        \gensync1/N174 ), .Q(\gensync1/N9 ) );
  INV3 U3304 ( .A(n1376), .Q(n874) );
  NOR21 U3305 ( .A(\gensync1/N176 ), .B(\gensync1/N177 ), .Q(n1376) );
  INV3 U3306 ( .A(reset_top), .Q(n653) );
  NOR21 U3307 ( .A(\gensync1/N180 ), .B(\gensync1/N179 ), .Q(\gensync1/n89 )
         );
  NOR21 U3308 ( .A(\gensync1/n102 ), .B(\gensync1/N74 ), .Q(\gensync1/N22 ) );
  BUF2 U3309 ( .A(\position1/N2452 ), .Q(n610) );
  BUF2 U3310 ( .A(\position1/N2460 ), .Q(n629) );
  BUF2 U3311 ( .A(\position1/N560 ), .Q(n516) );
  INV3 U3312 ( .A(reset_top), .Q(n652) );
  BUF2 U3313 ( .A(\position1/N2446 ), .Q(n598) );
  INV3 U3314 ( .A(reset_top), .Q(n651) );
  BUF2 U3315 ( .A(\position1/N2450 ), .Q(n606) );
  BUF2 U3316 ( .A(\position1/N2448 ), .Q(n602) );
  BUF2 U3317 ( .A(\position1/N2454 ), .Q(n616) );
  INV3 U3318 ( .A(\position1/n833 ), .Q(n691) );
  AOI221 U3319 ( .A(n484), .B(Y_barycentre_top[8]), .C(n634), .D(
        \position1/quot_y [8]), .Q(\position1/n833 ) );
  BUF2 U3320 ( .A(\position1/N2460 ), .Q(n632) );
  INV3 U3321 ( .A(\position1/n847 ), .Q(n678) );
  AOI221 U3322 ( .A(n484), .B(X_barycentre_top[4]), .C(n633), .D(
        \position1/quot_x [4]), .Q(\position1/n847 ) );
  INV3 U3323 ( .A(\position1/n838 ), .Q(n687) );
  AOI221 U3324 ( .A(n484), .B(Y_barycentre_top[4]), .C(n634), .D(
        \position1/quot_y [4]), .Q(\position1/n838 ) );
  INV3 U3325 ( .A(\position1/n835 ), .Q(n690) );
  AOI221 U3326 ( .A(n484), .B(Y_barycentre_top[7]), .C(n634), .D(
        \position1/quot_y [7]), .Q(\position1/n835 ) );
  INV3 U3327 ( .A(\position1/n836 ), .Q(n689) );
  AOI221 U3328 ( .A(n484), .B(Y_barycentre_top[6]), .C(n634), .D(
        \position1/quot_y [6]), .Q(\position1/n836 ) );
  INV3 U3329 ( .A(\position1/n846 ), .Q(n679) );
  AOI221 U3330 ( .A(n484), .B(X_barycentre_top[5]), .C(\position1/n834 ), .D(
        \position1/quot_x [5]), .Q(\position1/n846 ) );
  INV3 U3331 ( .A(\position1/n837 ), .Q(n688) );
  AOI221 U3332 ( .A(n484), .B(Y_barycentre_top[5]), .C(n634), .D(
        \position1/quot_y [5]), .Q(\position1/n837 ) );
  INV3 U3333 ( .A(\position1/n839 ), .Q(n686) );
  AOI221 U3334 ( .A(n484), .B(Y_barycentre_top[3]), .C(n634), .D(
        \position1/quot_y [3]), .Q(\position1/n839 ) );
  INV3 U3335 ( .A(\position1/n840 ), .Q(n685) );
  AOI221 U3336 ( .A(n484), .B(Y_barycentre_top[2]), .C(n634), .D(
        \position1/quot_y [2]), .Q(\position1/n840 ) );
  BUF2 U3337 ( .A(\position1/N2456 ), .Q(n619) );
  BUF2 U3338 ( .A(\position1/N2459 ), .Q(n626) );
  BUF2 U3339 ( .A(\position1/N2445 ), .Q(n593) );
  BUF2 U3340 ( .A(\position1/N560 ), .Q(n517) );
  INV3 U3341 ( .A(\image_process1/n62 ), .Q(n742) );
  NAND22 U3342 ( .A(reset_top), .B(b_top[7]), .Q(\image_process1/n62 ) );
  INV3 U3343 ( .A(\position1/n1183 ), .Q(n716) );
  NAND22 U3344 ( .A(b_out_proc[7]), .B(reset_top), .Q(\position1/n1183 ) );
  INV3 U3345 ( .A(\position1/n1192 ), .Q(n724) );
  NAND22 U3346 ( .A(g_out_proc[7]), .B(n649), .Q(\position1/n1192 ) );
  INV3 U3347 ( .A(\position1/n1193 ), .Q(n725) );
  NAND22 U3348 ( .A(g_out_proc[6]), .B(n649), .Q(\position1/n1193 ) );
  INV3 U3349 ( .A(\position1/n1194 ), .Q(n726) );
  NAND22 U3350 ( .A(g_out_proc[5]), .B(n649), .Q(\position1/n1194 ) );
  INV3 U3351 ( .A(\position1/n1195 ), .Q(n727) );
  NAND22 U3352 ( .A(g_out_proc[4]), .B(n649), .Q(\position1/n1195 ) );
  INV3 U3353 ( .A(\position1/n1184 ), .Q(n717) );
  NAND22 U3354 ( .A(b_out_proc[6]), .B(n649), .Q(\position1/n1184 ) );
  INV3 U3355 ( .A(\position1/n1185 ), .Q(n718) );
  NAND22 U3356 ( .A(b_out_proc[5]), .B(n649), .Q(\position1/n1185 ) );
  INV3 U3357 ( .A(\position1/n1186 ), .Q(n719) );
  NAND22 U3358 ( .A(b_out_proc[4]), .B(n649), .Q(\position1/n1186 ) );
  INV3 U3359 ( .A(\position1/n1188 ), .Q(n720) );
  NAND22 U3360 ( .A(b_out_proc[3]), .B(n649), .Q(\position1/n1188 ) );
  INV3 U3361 ( .A(\position1/n1189 ), .Q(n721) );
  NAND22 U3362 ( .A(b_out_proc[2]), .B(n649), .Q(\position1/n1189 ) );
  INV3 U3363 ( .A(\position1/n1190 ), .Q(n722) );
  NAND22 U3364 ( .A(b_out_proc[1]), .B(n649), .Q(\position1/n1190 ) );
  INV3 U3365 ( .A(\position1/n1191 ), .Q(n723) );
  NAND22 U3366 ( .A(b_out_proc[0]), .B(n649), .Q(\position1/n1191 ) );
  INV3 U3367 ( .A(\position1/n1200 ), .Q(n732) );
  NAND22 U3368 ( .A(r_out_proc[7]), .B(n649), .Q(\position1/n1200 ) );
  INV3 U3369 ( .A(\position1/n1201 ), .Q(n733) );
  NAND22 U3370 ( .A(r_out_proc[6]), .B(n649), .Q(\position1/n1201 ) );
  INV3 U3371 ( .A(\position1/n1202 ), .Q(n734) );
  NAND22 U3372 ( .A(r_out_proc[5]), .B(n649), .Q(\position1/n1202 ) );
  INV3 U3373 ( .A(\position1/n1203 ), .Q(n735) );
  NAND22 U3374 ( .A(r_out_proc[4]), .B(n649), .Q(\position1/n1203 ) );
  INV3 U3375 ( .A(\position1/n1204 ), .Q(n736) );
  NAND22 U3376 ( .A(r_out_proc[3]), .B(n649), .Q(\position1/n1204 ) );
  INV3 U3377 ( .A(\position1/n1205 ), .Q(n737) );
  NAND22 U3378 ( .A(r_out_proc[2]), .B(reset_top), .Q(\position1/n1205 ) );
  INV3 U3379 ( .A(\position1/n1206 ), .Q(n738) );
  NAND22 U3380 ( .A(r_out_proc[1]), .B(n649), .Q(\position1/n1206 ) );
  INV3 U3381 ( .A(\position1/n1207 ), .Q(n739) );
  NAND22 U3382 ( .A(r_out_proc[0]), .B(n649), .Q(\position1/n1207 ) );
  INV3 U3383 ( .A(\position1/n1196 ), .Q(n728) );
  NAND22 U3384 ( .A(g_out_proc[3]), .B(n649), .Q(\position1/n1196 ) );
  INV3 U3385 ( .A(\position1/n1197 ), .Q(n729) );
  NAND22 U3386 ( .A(g_out_proc[2]), .B(n649), .Q(\position1/n1197 ) );
  INV3 U3387 ( .A(\position1/n1198 ), .Q(n730) );
  NAND22 U3388 ( .A(g_out_proc[1]), .B(n649), .Q(\position1/n1198 ) );
  INV3 U3389 ( .A(\position1/n1199 ), .Q(n731) );
  NAND22 U3390 ( .A(g_out_proc[0]), .B(n649), .Q(\position1/n1199 ) );
  INV3 U3391 ( .A(\image_process1/n70 ), .Q(n750) );
  NAND22 U3392 ( .A(g_top[7]), .B(n648), .Q(\image_process1/n70 ) );
  INV3 U3393 ( .A(\image_process1/n71 ), .Q(n751) );
  NAND22 U3394 ( .A(g_top[6]), .B(n648), .Q(\image_process1/n71 ) );
  INV3 U3395 ( .A(\image_process1/n72 ), .Q(n752) );
  NAND22 U3396 ( .A(g_top[5]), .B(n648), .Q(\image_process1/n72 ) );
  INV3 U3397 ( .A(\image_process1/n73 ), .Q(n753) );
  NAND22 U3398 ( .A(g_top[4]), .B(n648), .Q(\image_process1/n73 ) );
  INV3 U3399 ( .A(\image_process1/n63 ), .Q(n743) );
  NAND22 U3400 ( .A(b_top[6]), .B(n648), .Q(\image_process1/n63 ) );
  INV3 U3401 ( .A(\image_process1/n64 ), .Q(n744) );
  NAND22 U3402 ( .A(b_top[5]), .B(n648), .Q(\image_process1/n64 ) );
  INV3 U3403 ( .A(\image_process1/n65 ), .Q(n745) );
  NAND22 U3404 ( .A(b_top[4]), .B(n648), .Q(\image_process1/n65 ) );
  INV3 U3405 ( .A(\image_process1/n66 ), .Q(n746) );
  NAND22 U3406 ( .A(b_top[3]), .B(n648), .Q(\image_process1/n66 ) );
  INV3 U3407 ( .A(\image_process1/n67 ), .Q(n747) );
  NAND22 U3408 ( .A(b_top[2]), .B(n648), .Q(\image_process1/n67 ) );
  INV3 U3409 ( .A(\image_process1/n68 ), .Q(n748) );
  NAND22 U3410 ( .A(b_top[1]), .B(n648), .Q(\image_process1/n68 ) );
  INV3 U3411 ( .A(\image_process1/n69 ), .Q(n749) );
  NAND22 U3412 ( .A(b_top[0]), .B(n648), .Q(\image_process1/n69 ) );
  INV3 U3413 ( .A(\image_process1/n78 ), .Q(n758) );
  NAND22 U3414 ( .A(r_top[7]), .B(reset_top), .Q(\image_process1/n78 ) );
  INV3 U3415 ( .A(\image_process1/n79 ), .Q(n759) );
  NAND22 U3416 ( .A(r_top[6]), .B(reset_top), .Q(\image_process1/n79 ) );
  INV3 U3417 ( .A(\image_process1/n80 ), .Q(n760) );
  NAND22 U3418 ( .A(r_top[5]), .B(reset_top), .Q(\image_process1/n80 ) );
  INV3 U3419 ( .A(\image_process1/n81 ), .Q(n761) );
  NAND22 U3420 ( .A(r_top[4]), .B(reset_top), .Q(\image_process1/n81 ) );
  INV3 U3421 ( .A(\image_process1/n82 ), .Q(n762) );
  NAND22 U3422 ( .A(r_top[3]), .B(reset_top), .Q(\image_process1/n82 ) );
  INV3 U3423 ( .A(\image_process1/n83 ), .Q(n763) );
  NAND22 U3424 ( .A(r_top[2]), .B(reset_top), .Q(\image_process1/n83 ) );
  INV3 U3425 ( .A(\image_process1/n84 ), .Q(n764) );
  NAND22 U3426 ( .A(r_top[1]), .B(reset_top), .Q(\image_process1/n84 ) );
  INV3 U3427 ( .A(\image_process1/n85 ), .Q(n765) );
  NAND22 U3428 ( .A(r_top[0]), .B(reset_top), .Q(\image_process1/n85 ) );
  INV3 U3429 ( .A(\image_process1/n74 ), .Q(n754) );
  NAND22 U3430 ( .A(g_top[3]), .B(reset_top), .Q(\image_process1/n74 ) );
  INV3 U3431 ( .A(\image_process1/n75 ), .Q(n755) );
  NAND22 U3432 ( .A(g_top[2]), .B(reset_top), .Q(\image_process1/n75 ) );
  INV3 U3433 ( .A(\image_process1/n76 ), .Q(n756) );
  NAND22 U3434 ( .A(g_top[1]), .B(reset_top), .Q(\image_process1/n76 ) );
  INV3 U3435 ( .A(\image_process1/n77 ), .Q(n757) );
  NAND22 U3436 ( .A(g_top[0]), .B(reset_top), .Q(\image_process1/n77 ) );
  NAND22 U3437 ( .A(\position1/x_sum [7]), .B(n519), .Q(\position1/n1571 ) );
  NAND22 U3438 ( .A(\position1/y_sum [7]), .B(n553), .Q(\position1/n1375 ) );
  NAND22 U3439 ( .A(\position1/N1529 ), .B(n519), .Q(\position1/n1570 ) );
  XNR21 U3440 ( .A(\position1/x_sum [8]), .B(n513), .Q(\position1/N1529 ) );
  NAND22 U3441 ( .A(\position1/N1946 ), .B(n553), .Q(\position1/n1374 ) );
  XNR21 U3442 ( .A(\position1/y_sum [8]), .B(n513), .Q(\position1/N1946 ) );
  NAND22 U3443 ( .A(\position1/N1533 ), .B(n519), .Q(\position1/n1566 ) );
  NAND22 U3444 ( .A(\position1/N1950 ), .B(n553), .Q(\position1/n1370 ) );
  NAND22 U3445 ( .A(\position1/N1535 ), .B(n518), .Q(\position1/n1564 ) );
  NAND22 U3446 ( .A(\position1/N1952 ), .B(n552), .Q(\position1/n1368 ) );
  NAND22 U3447 ( .A(\position1/N1537 ), .B(n518), .Q(\position1/n1562 ) );
  NAND22 U3448 ( .A(\position1/N1954 ), .B(n552), .Q(\position1/n1366 ) );
  NAND22 U3449 ( .A(\position1/N1539 ), .B(n518), .Q(\position1/n1560 ) );
  NAND22 U3450 ( .A(\position1/N1956 ), .B(n552), .Q(\position1/n1364 ) );
  NAND22 U3451 ( .A(\position1/N1541 ), .B(n518), .Q(\position1/n1558 ) );
  NAND22 U3452 ( .A(\position1/N1958 ), .B(n552), .Q(\position1/n1362 ) );
  NAND22 U3453 ( .A(\position1/N1543 ), .B(n518), .Q(\position1/n1556 ) );
  NAND22 U3454 ( .A(\position1/N1960 ), .B(n552), .Q(\position1/n1360 ) );
  NAND22 U3455 ( .A(\position1/N1531 ), .B(n519), .Q(\position1/n1568 ) );
  NAND22 U3456 ( .A(\position1/N1948 ), .B(n553), .Q(\position1/n1372 ) );
  NAND22 U3457 ( .A(\position1/N1545 ), .B(n518), .Q(\position1/n1554 ) );
  NAND22 U3458 ( .A(\position1/N1962 ), .B(n552), .Q(\position1/n1358 ) );
  AOI221 U3459 ( .A(\position1/x_sum [12]), .B(n248), .C(n2091), .D(n1340), 
        .Q(n2093) );
  INV3 U3460 ( .A(n2090), .Q(n1340) );
  AOI221 U3461 ( .A(n2089), .B(n1342), .C(n623), .D(n65), .Q(n2091) );
  NOR21 U3462 ( .A(n276), .B(\position1/x_sum [12]), .Q(n2090) );
  AOI221 U3463 ( .A(\position1/y_sum [12]), .B(n41), .C(n1757), .D(n1339), .Q(
        n1759) );
  INV3 U3464 ( .A(n1756), .Q(n1339) );
  AOI221 U3465 ( .A(n1755), .B(n1341), .C(n623), .D(n58), .Q(n1757) );
  NOR21 U3466 ( .A(n276), .B(\position1/y_sum [12]), .Q(n1756) );
  AOI221 U3467 ( .A(\position1/x_sum [14]), .B(n252), .C(n2095), .D(n1336), 
        .Q(n2097) );
  INV3 U3468 ( .A(n2094), .Q(n1336) );
  AOI221 U3469 ( .A(n2093), .B(n1338), .C(n620), .D(n64), .Q(n2095) );
  NOR21 U3470 ( .A(n45), .B(\position1/x_sum [14]), .Q(n2094) );
  AOI221 U3471 ( .A(\position1/y_sum [14]), .B(n280), .C(n1761), .D(n1335), 
        .Q(n1763) );
  INV3 U3472 ( .A(n1760), .Q(n1335) );
  AOI221 U3473 ( .A(n1759), .B(n1337), .C(n620), .D(n57), .Q(n1761) );
  NOR21 U3474 ( .A(n280), .B(\position1/y_sum [14]), .Q(n1760) );
  AOI221 U3475 ( .A(\position1/x_sum [16]), .B(n284), .C(n2099), .D(n1332), 
        .Q(n2101) );
  INV3 U3476 ( .A(n2098), .Q(n1332) );
  AOI221 U3477 ( .A(n2097), .B(n1334), .C(n616), .D(n63), .Q(n2099) );
  NOR21 U3478 ( .A(n284), .B(\position1/x_sum [16]), .Q(n2098) );
  AOI221 U3479 ( .A(\position1/y_sum [16]), .B(n256), .C(n1765), .D(n1331), 
        .Q(n1767) );
  INV3 U3480 ( .A(n1764), .Q(n1331) );
  AOI221 U3481 ( .A(n1763), .B(n1333), .C(n616), .D(n56), .Q(n1765) );
  NOR21 U3482 ( .A(n256), .B(\position1/y_sum [16]), .Q(n1764) );
  AOI221 U3483 ( .A(\position1/x_sum [18]), .B(n288), .C(n2103), .D(n1328), 
        .Q(n2105) );
  INV3 U3484 ( .A(n2102), .Q(n1328) );
  AOI221 U3485 ( .A(n2101), .B(n1330), .C(n611), .D(n62), .Q(n2103) );
  NOR21 U3486 ( .A(n46), .B(\position1/x_sum [18]), .Q(n2102) );
  AOI221 U3487 ( .A(\position1/y_sum [18]), .B(n259), .C(n1769), .D(n1327), 
        .Q(n1771) );
  INV3 U3488 ( .A(n1768), .Q(n1327) );
  AOI221 U3489 ( .A(n1767), .B(n1329), .C(n610), .D(n55), .Q(n1769) );
  NOR21 U3490 ( .A(n46), .B(\position1/y_sum [18]), .Q(n1768) );
  AOI221 U3491 ( .A(\position1/x_sum [20]), .B(n263), .C(n2107), .D(n1324), 
        .Q(n2109) );
  INV3 U3492 ( .A(n2106), .Q(n1324) );
  AOI221 U3493 ( .A(n2105), .B(n1326), .C(n606), .D(n61), .Q(n2107) );
  NOR21 U3494 ( .A(n43), .B(\position1/x_sum [20]), .Q(n2106) );
  AOI221 U3495 ( .A(\position1/y_sum [20]), .B(n292), .C(n1773), .D(n1323), 
        .Q(n1775) );
  INV3 U3496 ( .A(n1772), .Q(n1323) );
  AOI221 U3497 ( .A(n1771), .B(n1325), .C(n606), .D(n54), .Q(n1773) );
  NOR21 U3498 ( .A(n263), .B(\position1/y_sum [20]), .Q(n1772) );
  AOI221 U3499 ( .A(\position1/x_sum [22]), .B(n267), .C(n2111), .D(n1320), 
        .Q(n2113) );
  INV3 U3500 ( .A(n2110), .Q(n1320) );
  AOI221 U3501 ( .A(n2109), .B(n1322), .C(n602), .D(n60), .Q(n2111) );
  NOR21 U3502 ( .A(n42), .B(\position1/x_sum [22]), .Q(n2110) );
  AOI221 U3503 ( .A(\position1/y_sum [22]), .B(n267), .C(n1777), .D(n1319), 
        .Q(n1779) );
  INV3 U3504 ( .A(n1776), .Q(n1319) );
  AOI221 U3505 ( .A(n1775), .B(n1321), .C(n602), .D(n53), .Q(n1777) );
  NOR21 U3506 ( .A(n296), .B(\position1/y_sum [22]), .Q(n1776) );
  AOI221 U3507 ( .A(\position1/x_sum [10]), .B(n272), .C(n1344), .D(n2087), 
        .Q(n2089) );
  INV3 U3508 ( .A(n2086), .Q(n1344) );
  NAND22 U3509 ( .A(n630), .B(n51), .Q(n2087) );
  AOI221 U3510 ( .A(\position1/y_sum [10]), .B(n245), .C(n1343), .D(n1753), 
        .Q(n1755) );
  INV3 U3511 ( .A(n1752), .Q(n1343) );
  NAND22 U3512 ( .A(n631), .B(n50), .Q(n1753) );
  NOR40 U3513 ( .A(\position1/x_sum [7]), .B(\position1/x_sum [6]), .C(
        \position1/x_sum [5]), .D(\position1/x_sum [4]), .Q(n2081) );
  NOR40 U3514 ( .A(\position1/y_sum [7]), .B(\position1/y_sum [6]), .C(
        \position1/y_sum [5]), .D(\position1/y_sum [4]), .Q(n1747) );
  NAND22 U3515 ( .A(\position1/x_sum [4]), .B(n519), .Q(\position1/n1574 ) );
  NAND22 U3516 ( .A(\position1/y_sum [4]), .B(n553), .Q(\position1/n1378 ) );
  NAND22 U3517 ( .A(\position1/x_sum [3]), .B(n519), .Q(\position1/n1575 ) );
  NAND22 U3518 ( .A(\position1/y_sum [3]), .B(n553), .Q(\position1/n1379 ) );
  NAND22 U3519 ( .A(\position1/x_sum [5]), .B(n519), .Q(\position1/n1573 ) );
  NAND22 U3520 ( .A(\position1/y_sum [5]), .B(n553), .Q(\position1/n1377 ) );
  NAND22 U3521 ( .A(\position1/x_sum [6]), .B(n519), .Q(\position1/n1572 ) );
  NAND22 U3522 ( .A(\position1/y_sum [6]), .B(n553), .Q(\position1/n1376 ) );
  NAND22 U3523 ( .A(\position1/N1521 ), .B(n519), .Q(\position1/n1578 ) );
  NAND22 U3524 ( .A(\position1/N1938 ), .B(n553), .Q(\position1/n1382 ) );
  NAND22 U3525 ( .A(\position1/x_sum [1]), .B(n520), .Q(\position1/n1577 ) );
  NAND22 U3526 ( .A(\position1/y_sum [1]), .B(n554), .Q(\position1/n1381 ) );
  NAND22 U3527 ( .A(\position1/x_sum [2]), .B(n519), .Q(\position1/n1576 ) );
  NAND22 U3528 ( .A(\position1/y_sum [2]), .B(n553), .Q(\position1/n1380 ) );
  NOR21 U3529 ( .A(n586), .B(n2116), .Q(\position1/N1519 ) );
  AOI221 U3530 ( .A(\position1/x_sum [24]), .B(n300), .C(n2115), .D(n1346), 
        .Q(n2116) );
  INV3 U3531 ( .A(n2114), .Q(n1346) );
  AOI221 U3532 ( .A(n2113), .B(n1318), .C(n598), .D(n59), .Q(n2115) );
  NOR21 U3533 ( .A(n586), .B(n1782), .Q(\position1/N1936 ) );
  AOI221 U3534 ( .A(\position1/y_sum [24]), .B(n300), .C(n1781), .D(n1345), 
        .Q(n1782) );
  INV3 U3535 ( .A(n1780), .Q(n1345) );
  AOI221 U3536 ( .A(n1779), .B(n1099), .C(n598), .D(n52), .Q(n1781) );
  NOR21 U3537 ( .A(n300), .B(\position1/x_sum [24]), .Q(n2114) );
  NOR21 U3538 ( .A(n300), .B(\position1/y_sum [24]), .Q(n1780) );
  INV3 U3539 ( .A(n2083), .Q(n1348) );
  AOI221 U3540 ( .A(n2082), .B(n2081), .C(n516), .D(n49), .Q(n2083) );
  NOR40 U3541 ( .A(\position1/x_sum [3]), .B(\position1/x_sum [2]), .C(
        \position1/x_sum [1]), .D(\position1/N1521 ), .Q(n2082) );
  INV3 U3542 ( .A(n1749), .Q(n1347) );
  AOI221 U3543 ( .A(n1748), .B(n1747), .C(n516), .D(n48), .Q(n1749) );
  NOR40 U3544 ( .A(\position1/y_sum [3]), .B(\position1/y_sum [2]), .C(
        \position1/y_sum [1]), .D(\position1/N1938 ), .Q(n1748) );
  INV3 U3545 ( .A(n165), .Q(\position1/sub_216/carry [9]) );
  NOR21 U3546 ( .A(n513), .B(\position1/x_sum [8]), .Q(n165) );
  INV3 U3547 ( .A(n164), .Q(\position1/sub_226/carry [9]) );
  NOR21 U3548 ( .A(n513), .B(\position1/y_sum [8]), .Q(n164) );
  BUF2 U3549 ( .A(\position1/N2452 ), .Q(n609) );
  BUF2 U3550 ( .A(\position1/N2445 ), .Q(n591) );
  BUF2 U3551 ( .A(\position1/N2459 ), .Q(n624) );
  BUF2 U3552 ( .A(\position1/N2456 ), .Q(n617) );
  BUF2 U3553 ( .A(\position1/N2450 ), .Q(n603) );
  BUF2 U3554 ( .A(\position1/N2448 ), .Q(n599) );
  BUF2 U3555 ( .A(\position1/N2458 ), .Q(n622) );
  BUF2 U3556 ( .A(\position1/N2446 ), .Q(n595) );
  BUF2 U3557 ( .A(\position1/N2454 ), .Q(n612) );
  BUF2 U3558 ( .A(\position1/N2454 ), .Q(n614) );
  BUF2 U3559 ( .A(\position1/N2452 ), .Q(n611) );
  LOGIC1 U3560 ( .Q(\position1/n283 ) );
  LOGIC0 U3561 ( .Q(\*Logic0* ) );
  OAI212 U3562 ( .A(n1368), .B(n1367), .C(n1366), .Q(n1369) );
  OAI212 U3563 ( .A(\gensync1/N181 ), .B(\gensync1/N182 ), .C(\gensync1/N180 ), 
        .Q(n1378) );
  OAI212 U3564 ( .A(\gensync1/N181 ), .B(\gensync1/N182 ), .C(\gensync1/N180 ), 
        .Q(n1380) );
  OAI212 U3565 ( .A(n1384), .B(n5), .C(n33), .Q(n1385) );
  OAI212 U3566 ( .A(Y_barycentre_top[3]), .B(n801), .C(n1392), .Q(n1393) );
  OAI212 U3567 ( .A(\position1/N2407 ), .B(n24), .C(n1393), .Q(n1394) );
  OAI222 U3568 ( .A(n1395), .B(n1394), .C(Y_barycentre_top[4]), .D(n797), .Q(
        n1396) );
  OAI222 U3569 ( .A(\position1/N2409 ), .B(n28), .C(n1397), .D(n1396), .Q(
        n1398) );
  OAI222 U3570 ( .A(n1399), .B(n1398), .C(Y_barycentre_top[6]), .D(n789), .Q(
        n1400) );
  OAI222 U3571 ( .A(\position1/N2411 ), .B(n32), .C(n1401), .D(n1400), .Q(
        n1402) );
  OAI222 U3572 ( .A(n1403), .B(n1402), .C(Y_barycentre_top[8]), .D(n779), .Q(
        \position1/N2413 ) );
  OAI212 U3573 ( .A(X_barycentre_top[3]), .B(n841), .C(n1407), .Q(n1408) );
  OAI212 U3574 ( .A(\position1/N2396 ), .B(n19), .C(n1408), .Q(n1409) );
  OAI222 U3575 ( .A(n1410), .B(n1409), .C(X_barycentre_top[4]), .D(n840), .Q(
        n1411) );
  OAI222 U3576 ( .A(\position1/N2398 ), .B(n22), .C(n1412), .D(n1411), .Q(
        n1413) );
  OAI222 U3577 ( .A(n1414), .B(n1413), .C(X_barycentre_top[6]), .D(n838), .Q(
        n1415) );
  OAI222 U3578 ( .A(\position1/N2400 ), .B(n27), .C(n1416), .D(n1415), .Q(
        n1417) );
  OAI222 U3579 ( .A(n1418), .B(n1417), .C(X_barycentre_top[8]), .D(n836), .Q(
        \position1/N2402 ) );
  OAI212 U3580 ( .A(\position1/N2385 ), .B(n24), .C(n1422), .Q(n1423) );
  OAI212 U3581 ( .A(Y_barycentre_top[3]), .B(n802), .C(n1423), .Q(n1424) );
  OAI222 U3582 ( .A(n1425), .B(n1424), .C(\position1/N2386 ), .D(n26), .Q(
        n1426) );
  OAI222 U3583 ( .A(Y_barycentre_top[5]), .B(n794), .C(n1427), .D(n1426), .Q(
        n1428) );
  OAI222 U3584 ( .A(n1429), .B(n1428), .C(\position1/N2388 ), .D(n31), .Q(
        n1430) );
  OAI222 U3585 ( .A(Y_barycentre_top[7]), .B(n786), .C(n1431), .D(n1430), .Q(
        n1432) );
  OAI222 U3586 ( .A(n1433), .B(n1432), .C(\position1/N2390 ), .D(n30), .Q(
        \position1/N2391 ) );
  OAI212 U3587 ( .A(\position1/N2375 ), .B(n19), .C(n1437), .Q(n1438) );
  OAI212 U3588 ( .A(X_barycentre_top[3]), .B(n849), .C(n1438), .Q(n1439) );
  OAI222 U3589 ( .A(n1440), .B(n1439), .C(\position1/N2376 ), .D(n20), .Q(
        n1441) );
  OAI222 U3590 ( .A(X_barycentre_top[5]), .B(n847), .C(n1442), .D(n1441), .Q(
        n1443) );
  OAI222 U3591 ( .A(n1444), .B(n1443), .C(\position1/N2378 ), .D(n25), .Q(
        n1445) );
  OAI222 U3592 ( .A(X_barycentre_top[7]), .B(n845), .C(n1446), .D(n1445), .Q(
        n1447) );
  OAI222 U3593 ( .A(n1448), .B(n1447), .C(\position1/N2380 ), .D(n29), .Q(
        \position1/N2381 ) );
  OAI212 U3594 ( .A(n1450), .B(n629), .C(\position1/n1231 ), .Q(n1449) );
  OAI222 U3595 ( .A(\position1/n1224 ), .B(n471), .C(n895), .D(n894), .Q(n1466) );
  OAI222 U3596 ( .A(n1466), .B(n1465), .C(n259), .D(n893), .Q(n1467) );
  OAI212 U3597 ( .A(n593), .B(\position1/n1264 ), .C(n1555), .Q(n1557) );
  OAI222 U3598 ( .A(n1564), .B(n1563), .C(n515), .D(\position1/n1304 ), .Q(
        n1565) );
  OAI222 U3599 ( .A(n988), .B(n628), .C(n1566), .D(n1565), .Q(n1567) );
  OAI222 U3600 ( .A(n1568), .B(n1567), .C(n624), .D(\position1/n1302 ), .Q(
        n1569) );
  OAI222 U3601 ( .A(n986), .B(n37), .C(n1570), .D(n1569), .Q(n1571) );
  OAI222 U3602 ( .A(n1572), .B(n1571), .C(n468), .D(\position1/n1300 ), .Q(
        n1573) );
  OAI222 U3603 ( .A(n984), .B(n47), .C(n1574), .D(n1573), .Q(n1575) );
  OAI222 U3604 ( .A(n1576), .B(n1575), .C(n469), .D(\position1/n1298 ), .Q(
        n1577) );
  OAI222 U3605 ( .A(n982), .B(n254), .C(n1578), .D(n1577), .Q(n1579) );
  OAI222 U3606 ( .A(n1580), .B(n1579), .C(n471), .D(\position1/n1296 ), .Q(
        n1581) );
  OAI222 U3607 ( .A(n980), .B(n286), .C(n1582), .D(n1581), .Q(n1583) );
  OAI222 U3608 ( .A(n1584), .B(n1583), .C(n473), .D(\position1/n1294 ), .Q(
        n1585) );
  OAI222 U3609 ( .A(n978), .B(n38), .C(n1586), .D(n1585), .Q(n1587) );
  OAI222 U3610 ( .A(n1588), .B(n1587), .C(n474), .D(\position1/n1292 ), .Q(
        n1589) );
  OAI222 U3611 ( .A(n976), .B(n39), .C(n1590), .D(n1589), .Q(n1591) );
  OAI222 U3612 ( .A(n1592), .B(n1591), .C(n475), .D(\position1/n1290 ), .Q(
        n1593) );
  OAI222 U3613 ( .A(n1604), .B(n1019), .C(n515), .D(\position1/n1328 ), .Q(
        n1605) );
  OAI222 U3614 ( .A(n1018), .B(n628), .C(n1017), .D(n1605), .Q(n1606) );
  OAI222 U3615 ( .A(n1015), .B(n1606), .C(n626), .D(\position1/n1326 ), .Q(
        n1607) );
  OAI222 U3616 ( .A(n1014), .B(n37), .C(n1013), .D(n1607), .Q(n1608) );
  OAI222 U3617 ( .A(n1011), .B(n1608), .C(\position1/N2457 ), .D(
        \position1/n1324 ), .Q(n1609) );
  OAI222 U3618 ( .A(n1009), .B(n252), .C(n1610), .D(n1609), .Q(n1611) );
  OAI212 U3619 ( .A(n631), .B(n1044), .C(n1639), .Q(n1640) );
  OAI212 U3620 ( .A(\position1/N2073 ), .B(n628), .C(n1640), .Q(n1641) );
  OAI222 U3621 ( .A(n1642), .B(n1641), .C(n626), .D(n1043), .Q(n1643) );
  OAI222 U3622 ( .A(\position1/N2075 ), .B(n37), .C(n1644), .D(n1643), .Q(
        n1645) );
  OAI222 U3623 ( .A(n1646), .B(n1645), .C(n468), .D(n1041), .Q(n1647) );
  OAI222 U3624 ( .A(\position1/N2077 ), .B(n47), .C(n1648), .D(n1647), .Q(
        n1649) );
  OAI222 U3625 ( .A(n1650), .B(n1649), .C(n470), .D(n1039), .Q(n1651) );
  OAI222 U3626 ( .A(\position1/N2079 ), .B(n282), .C(n1652), .D(n1651), .Q(
        n1653) );
  OAI222 U3627 ( .A(n1654), .B(n1653), .C(\position1/N2453 ), .D(n1037), .Q(
        n1655) );
  OAI222 U3628 ( .A(\position1/N2081 ), .B(n286), .C(n1656), .D(n1655), .Q(
        n1657) );
  OAI222 U3629 ( .A(n1658), .B(n1657), .C(n473), .D(n1035), .Q(n1659) );
  OAI222 U3630 ( .A(\position1/N2083 ), .B(n38), .C(n1660), .D(n1659), .Q(
        n1661) );
  OAI222 U3631 ( .A(n1662), .B(n1661), .C(\position1/N2449 ), .D(n1033), .Q(
        n1663) );
  OAI222 U3632 ( .A(\position1/N2085 ), .B(n39), .C(n1664), .D(n1663), .Q(
        n1665) );
  OAI222 U3633 ( .A(n1666), .B(n1665), .C(\position1/N2447 ), .D(n1031), .Q(
        n1667) );
  OAI222 U3634 ( .A(\position1/N2087 ), .B(n67), .C(n1668), .D(n1667), .Q(
        n1669) );
  OAI222 U3635 ( .A(n1670), .B(n1669), .C(n593), .D(n1028), .Q(n1671) );
  OAI212 U3636 ( .A(n1671), .B(n588), .C(\position1/N2089 ), .Q(n1673) );
  OAI212 U3637 ( .A(n631), .B(\position1/n1350 ), .C(n1678), .Q(n1679) );
  OAI212 U3638 ( .A(n1079), .B(n628), .C(n1679), .Q(n1680) );
  OAI222 U3639 ( .A(n1076), .B(n1680), .C(n626), .D(\position1/n1349 ), .Q(
        n1681) );
  OAI222 U3640 ( .A(n1072), .B(n276), .C(n1682), .D(n1681), .Q(n1683) );
  IMAJ31 U3641 ( .A(n1081), .B(n586), .C(n1746), .Q(\position1/N1988 ) );
  OAI212 U3642 ( .A(n48), .B(n515), .C(n1347), .Q(n1751) );
  OAI222 U3643 ( .A(n1751), .B(n1750), .C(n272), .D(\position1/y_sum [10]), 
        .Q(n1752) );
  OAI212 U3644 ( .A(n1784), .B(n631), .C(\position1/n1427 ), .Q(n1783) );
  OAI222 U3645 ( .A(\position1/n1420 ), .B(\position1/N2453 ), .C(n1114), .D(
        n1113), .Q(n1800) );
  OAI222 U3646 ( .A(n1800), .B(n1799), .C(n259), .D(n1112), .Q(n1801) );
  OAI212 U3647 ( .A(n594), .B(\position1/n1460 ), .C(n1889), .Q(n1891) );
  OAI222 U3648 ( .A(n1898), .B(n1897), .C(n516), .D(\position1/n1500 ), .Q(
        n1899) );
  OAI222 U3649 ( .A(n1207), .B(n628), .C(n1900), .D(n1899), .Q(n1901) );
  OAI222 U3650 ( .A(n1902), .B(n1901), .C(n626), .D(\position1/n1498 ), .Q(
        n1903) );
  OAI222 U3651 ( .A(n1205), .B(n37), .C(n1904), .D(n1903), .Q(n1905) );
  OAI222 U3652 ( .A(n1906), .B(n1905), .C(\position1/N2457 ), .D(
        \position1/n1496 ), .Q(n1907) );
  OAI222 U3653 ( .A(n1203), .B(n47), .C(n1908), .D(n1907), .Q(n1909) );
  OAI222 U3654 ( .A(n1910), .B(n1909), .C(n469), .D(\position1/n1494 ), .Q(
        n1911) );
  OAI222 U3655 ( .A(n1201), .B(n254), .C(n1912), .D(n1911), .Q(n1913) );
  OAI222 U3656 ( .A(n1914), .B(n1913), .C(n471), .D(\position1/n1492 ), .Q(
        n1915) );
  OAI222 U3657 ( .A(n1199), .B(n286), .C(n1916), .D(n1915), .Q(n1917) );
  OAI222 U3658 ( .A(n1918), .B(n1917), .C(n473), .D(\position1/n1490 ), .Q(
        n1919) );
  OAI222 U3659 ( .A(n1197), .B(n38), .C(n1920), .D(n1919), .Q(n1921) );
  OAI222 U3660 ( .A(n1922), .B(n1921), .C(n474), .D(\position1/n1488 ), .Q(
        n1923) );
  OAI222 U3661 ( .A(n1195), .B(n39), .C(n1924), .D(n1923), .Q(n1925) );
  OAI222 U3662 ( .A(n1926), .B(n1925), .C(n475), .D(\position1/n1486 ), .Q(
        n1927) );
  OAI222 U3663 ( .A(n1938), .B(n1238), .C(n516), .D(\position1/n1524 ), .Q(
        n1939) );
  OAI222 U3664 ( .A(n1237), .B(n628), .C(n1236), .D(n1939), .Q(n1940) );
  OAI222 U3665 ( .A(n1234), .B(n1940), .C(n626), .D(\position1/n1522 ), .Q(
        n1941) );
  OAI222 U3666 ( .A(n1233), .B(n37), .C(n1232), .D(n1941), .Q(n1942) );
  OAI222 U3667 ( .A(n1230), .B(n1942), .C(n468), .D(\position1/n1520 ), .Q(
        n1943) );
  OAI222 U3668 ( .A(n1228), .B(n45), .C(n1944), .D(n1943), .Q(n1945) );
  OAI212 U3669 ( .A(n631), .B(n1263), .C(n1973), .Q(n1974) );
  OAI212 U3670 ( .A(\position1/N1656 ), .B(n628), .C(n1974), .Q(n1975) );
  OAI222 U3671 ( .A(n1976), .B(n1975), .C(n626), .D(n1262), .Q(n1977) );
  OAI222 U3672 ( .A(\position1/N1658 ), .B(n37), .C(n1978), .D(n1977), .Q(
        n1979) );
  OAI222 U3673 ( .A(n1980), .B(n1979), .C(\position1/N2457 ), .D(n1260), .Q(
        n1981) );
  OAI222 U3674 ( .A(\position1/N1660 ), .B(n47), .C(n1982), .D(n1981), .Q(
        n1983) );
  OAI222 U3675 ( .A(n1984), .B(n1983), .C(n470), .D(n1258), .Q(n1985) );
  OAI222 U3676 ( .A(\position1/N1662 ), .B(n100), .C(n1986), .D(n1985), .Q(
        n1987) );
  OAI222 U3677 ( .A(n1988), .B(n1987), .C(\position1/N2453 ), .D(n1256), .Q(
        n1989) );
  OAI222 U3678 ( .A(\position1/N1664 ), .B(n286), .C(n1990), .D(n1989), .Q(
        n1991) );
  OAI222 U3679 ( .A(n1992), .B(n1991), .C(n473), .D(n1254), .Q(n1993) );
  OAI222 U3680 ( .A(\position1/N1666 ), .B(n38), .C(n1994), .D(n1993), .Q(
        n1995) );
  OAI222 U3681 ( .A(n1996), .B(n1995), .C(\position1/N2449 ), .D(n1252), .Q(
        n1997) );
  OAI222 U3682 ( .A(\position1/N1668 ), .B(n39), .C(n1998), .D(n1997), .Q(
        n1999) );
  OAI222 U3683 ( .A(n2000), .B(n1999), .C(\position1/N2447 ), .D(n1250), .Q(
        n2001) );
  OAI222 U3684 ( .A(\position1/N1670 ), .B(n67), .C(n2002), .D(n2001), .Q(
        n2003) );
  OAI222 U3685 ( .A(n2004), .B(n2003), .C(n593), .D(n1247), .Q(n2005) );
  OAI212 U3686 ( .A(n2005), .B(n589), .C(\position1/N1672 ), .Q(n2007) );
  OAI212 U3687 ( .A(n631), .B(\position1/n1546 ), .C(n2012), .Q(n2013) );
  OAI212 U3688 ( .A(n1298), .B(n628), .C(n2013), .Q(n2014) );
  OAI222 U3689 ( .A(n1295), .B(n2014), .C(n626), .D(\position1/n1545 ), .Q(
        n2015) );
  OAI222 U3690 ( .A(n1291), .B(n248), .C(n2016), .D(n2015), .Q(n2017) );
  IMAJ31 U3691 ( .A(n1300), .B(n586), .C(n2080), .Q(\position1/N1571 ) );
  OAI212 U3692 ( .A(n49), .B(n515), .C(n1348), .Q(n2085) );
  OAI222 U3693 ( .A(n2085), .B(n2084), .C(n66), .D(\position1/x_sum [10]), .Q(
        n2086) );
  OAI212 U3694 ( .A(n2119), .B(n2118), .C(n2117), .Q(n2120) );
endmodule

