../../BENCH/bench_position.vhd