../../VHD/constants.vhd