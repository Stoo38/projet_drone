../../BENCH/test_div.vhd