
module top_ppm ( i_clk_top, i_reset_n_top, i_sel_top, o_ppm_top );
  input [1:0] i_sel_top;
  input i_clk_top, i_reset_n_top;
  output o_ppm_top;
  wire   \send_ppm1/n95 , \send_ppm1/n94 , \send_ppm1/n93 , \send_ppm1/n92 ,
         \send_ppm1/n91 , \send_ppm1/n90 , \send_ppm1/n89 , \send_ppm1/n88 ,
         \send_ppm1/n87 , \send_ppm1/n86 , \send_ppm1/n85 , \send_ppm1/n84 ,
         \send_ppm1/n83 , \send_ppm1/n82 , \send_ppm1/n81 , \send_ppm1/n80 ,
         \send_ppm1/n79 , \send_ppm1/n78 , \send_ppm1/n77 , \send_ppm1/n76 ,
         \send_ppm1/n75 , \send_ppm1/n74 , \send_ppm1/n73 , \send_ppm1/n72 ,
         \send_ppm1/n71 , \send_ppm1/n70 , \send_ppm1/n69 , \send_ppm1/n68 ,
         \send_ppm1/n67 , \send_ppm1/n66 , \send_ppm1/n65 , \send_ppm1/n64 ,
         \send_ppm1/n63 , \send_ppm1/n62 , \send_ppm1/n61 , \send_ppm1/n60 ,
         \send_ppm1/n59 , \send_ppm1/n58 , \send_ppm1/n57 , \send_ppm1/n55 ,
         \send_ppm1/n53 , \send_ppm1/dp_cluster_4/N218 ,
         \send_ppm1/dp_cluster_4/N219 , \send_ppm1/dp_cluster_4/N220 ,
         \send_ppm1/dp_cluster_4/N221 , \send_ppm1/dp_cluster_4/N223 ,
         \send_ppm1/dp_cluster_3/N233 , \send_ppm1/dp_cluster_3/N234 ,
         \send_ppm1/dp_cluster_3/N235 , \send_ppm1/dp_cluster_3/N236 ,
         \send_ppm1/dp_cluster_3/N238 , \send_ppm1/dp_cluster_2/N248 ,
         \send_ppm1/dp_cluster_2/N249 , \send_ppm1/dp_cluster_2/N250 ,
         \send_ppm1/dp_cluster_2/N251 , \send_ppm1/dp_cluster_2/N253 ,
         \send_ppm1/dp_cluster_1/N263 , \send_ppm1/dp_cluster_1/N264 ,
         \send_ppm1/dp_cluster_1/N265 , \send_ppm1/dp_cluster_1/N266 ,
         \send_ppm1/dp_cluster_1/N268 , \send_ppm1/dp_cluster_0/N18 ,
         \send_ppm1/dp_cluster_0/N19 , \send_ppm1/dp_cluster_0/N20 ,
         \send_ppm1/dp_cluster_0/N21 , \send_ppm1/dp_cluster_0/N22 ,
         \send_ppm1/dp_cluster_0/N23 , \send_ppm1/dp_cluster_0/N24 ,
         \send_ppm1/dp_cluster_0/N25 , \send_ppm1/dp_cluster_0/N26 ,
         \send_ppm1/dp_cluster_0/N27 , \send_ppm1/dp_cluster_0/N278 ,
         \send_ppm1/dp_cluster_0/N279 , \send_ppm1/dp_cluster_0/N28 ,
         \send_ppm1/dp_cluster_0/N280 , \send_ppm1/dp_cluster_0/N281 ,
         \send_ppm1/dp_cluster_0/N282 , \send_ppm1/dp_cluster_0/N283 ,
         \send_ppm1/dp_cluster_0/N284 , \send_ppm1/dp_cluster_0/N285 ,
         \send_ppm1/dp_cluster_0/N286 , \send_ppm1/dp_cluster_0/N287 ,
         \send_ppm1/dp_cluster_0/N288 , \send_ppm1/dp_cluster_0/N289 ,
         \send_ppm1/dp_cluster_0/N29 , \send_ppm1/dp_cluster_0/N290 ,
         \send_ppm1/dp_cluster_0/N291 , \send_ppm1/dp_cluster_0/N292 ,
         \send_ppm1/dp_cluster_0/N293 , \send_ppm1/dp_cluster_0/N294 ,
         \send_ppm1/dp_cluster_0/N295 , \send_ppm1/dp_cluster_0/N296 ,
         \send_ppm1/dp_cluster_0/N30 , \send_ppm1/dp_cluster_0/N31 ,
         \send_ppm1/dp_cluster_0/N38 , \send_ppm1/dp_cluster_0/N39 ,
         \send_ppm1/dp_cluster_0/N40 , \send_ppm1/dp_cluster_0/N41 ,
         \send_ppm1/dp_cluster_0/N42 , \send_ppm1/dp_cluster_0/N43 ,
         \send_ppm1/dp_cluster_0/N44 , \send_ppm1/dp_cluster_0/N45 ,
         \send_ppm1/dp_cluster_0/N46 , \send_ppm1/dp_cluster_0/N47 ,
         \send_ppm1/dp_cluster_0/N48 , \send_ppm1/dp_cluster_0/N49 ,
         \send_ppm1/dp_cluster_0/N50 , \send_ppm1/dp_cluster_0/N51 ,
         \send_ppm1/N198 , \send_ppm1/N197 , \send_ppm1/N196 ,
         \send_ppm1/N195 , \send_ppm1/N194 , \send_ppm1/N193 ,
         \send_ppm1/N192 , \send_ppm1/N191 , \send_ppm1/N190 ,
         \send_ppm1/N189 , \send_ppm1/N188 , \send_ppm1/N187 ,
         \send_ppm1/N186 , \send_ppm1/N185 , \send_ppm1/N184 ,
         \send_ppm1/N183 , \send_ppm1/N182 , \send_ppm1/N181 ,
         \send_ppm1/N180 , \send_ppm1/N179 , \send_ppm1/N169 ,
         \send_ppm1/N163 , \send_ppm1/N156 , \send_ppm1/N148 , \send_ppm1/N82 ,
         \send_ppm1/N81 , \send_ppm1/sig_in_init ,
         \send_ppm1/local_counter1/n22 , \send_ppm1/local_counter1/N65 ,
         \send_ppm1/local_counter1/N64 , \send_ppm1/local_counter1/N63 ,
         \send_ppm1/local_counter1/N62 , \send_ppm1/local_counter1/N61 ,
         \send_ppm1/local_counter1/N60 , \send_ppm1/local_counter1/N59 ,
         \send_ppm1/local_counter1/N58 , \send_ppm1/local_counter1/N57 ,
         \send_ppm1/local_counter1/N56 , \send_ppm1/local_counter1/N55 ,
         \send_ppm1/local_counter1/N54 , \send_ppm1/local_counter1/N53 ,
         \send_ppm1/local_counter1/N52 , \send_ppm1/local_counter1/N51 ,
         \send_ppm1/local_counter1/N50 , \send_ppm1/local_counter1/N49 ,
         \send_ppm1/local_counter1/N48 , \send_ppm1/local_counter1/N47 ,
         \send_ppm1/local_counter1/N46 , \send_ppm1/local_counter1/N24 ,
         \send_ppm1/local_counter1/N23 , \send_ppm1/local_counter1/N22 ,
         \send_ppm1/local_counter1/N21 , \send_ppm1/local_counter1/N20 ,
         \send_ppm1/local_counter1/N19 , \send_ppm1/local_counter1/N18 ,
         \send_ppm1/local_counter1/N17 , \send_ppm1/local_counter1/N16 ,
         \send_ppm1/local_counter1/N15 , \send_ppm1/local_counter1/N14 ,
         \send_ppm1/local_counter1/N13 , \send_ppm1/local_counter1/N12 ,
         \send_ppm1/local_counter1/N11 , \send_ppm1/local_counter1/N10 ,
         \send_ppm1/local_counter1/N9 , \send_ppm1/local_counter1/N8 ,
         \send_ppm1/local_counter1/N7 ,
         \send_ppm1/dp_cluster_1/mult_114/A2[8] ,
         \send_ppm1/dp_cluster_1/mult_114/A2[12] ,
         \send_ppm1/dp_cluster_1/mult_114/A1[11] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[1][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[2][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[3][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[4][1] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[4][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[5][1] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[5][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[6][1] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[6][5] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[7][1] ,
         \send_ppm1/dp_cluster_1/mult_114/SUMB[7][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[1][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[2][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[3][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][1] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][1] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][1] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][5] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][1] ,
         \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][5] ,
         \send_ppm1/dp_cluster_2/mult_117/A2[8] ,
         \send_ppm1/dp_cluster_2/mult_117/A2[12] ,
         \send_ppm1/dp_cluster_2/mult_117/A1[11] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[1][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[2][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[3][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[4][1] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[4][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[5][1] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[5][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[6][1] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[6][5] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[7][1] ,
         \send_ppm1/dp_cluster_2/mult_117/SUMB[7][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[1][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[2][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[3][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][1] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][1] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][1] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][5] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][1] ,
         \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][5] ,
         \send_ppm1/dp_cluster_3/mult_120/A2[8] ,
         \send_ppm1/dp_cluster_3/mult_120/A2[12] ,
         \send_ppm1/dp_cluster_3/mult_120/A1[11] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[1][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[2][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[3][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[4][1] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[4][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[5][1] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[5][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[6][1] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[6][5] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[7][1] ,
         \send_ppm1/dp_cluster_3/mult_120/SUMB[7][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[1][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[2][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[3][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][1] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][1] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][1] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][5] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][1] ,
         \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][5] ,
         \send_ppm1/dp_cluster_4/mult_123/A2[8] ,
         \send_ppm1/dp_cluster_4/mult_123/A2[12] ,
         \send_ppm1/dp_cluster_4/mult_123/A1[11] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[1][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[2][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[3][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[4][1] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[4][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[5][1] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[5][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[6][1] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[6][5] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[7][1] ,
         \send_ppm1/dp_cluster_4/mult_123/SUMB[7][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[1][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[2][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[3][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][1] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][1] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][1] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][5] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][1] ,
         \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][5] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363;
  wire   [31:0] sig_reg;
  wire   [2:0] \send_ppm1/sig_state ;
  wire   [2:0] \send_ppm1/current_state ;
  wire   [15:0] \send_ppm1/sig_cyclesTrame4 ;
  wire   [15:0] \send_ppm1/sig_cyclesTrame3 ;
  wire   [15:0] \send_ppm1/sig_cyclesTrame2 ;
  wire   [15:0] \send_ppm1/sig_cyclesTrame1 ;
  wire   [31:0] \send_ppm1/sig_reg_storage ;
  wire   [19:0] \send_ppm1/sig_out_local_count ;
  wire   [19:0] \send_ppm1/local_counter1/v_val ;
  wire   [19:2] \send_ppm1/local_counter1/add_34/carry ;
  wire   [20:0] \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry ;
  wire   [19:1] \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry ;
  wire   [19:1] \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry ;
  wire   [20:0] \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry ;
  wire   [16:1] \send_ppm1/dp_cluster_1/sub_114_cf/carry ;
  wire   [16:1] \send_ppm1/dp_cluster_2/sub_117_cf/carry ;
  wire   [16:1] \send_ppm1/dp_cluster_3/sub_120_cf/carry ;
  wire   [16:1] \send_ppm1/dp_cluster_4/sub_123_cf/carry ;
  assign sig_reg[31] = i_sel_top[1];
  assign sig_reg[30] = i_sel_top[0];

  OAI222 \send_ppm1/U39  ( .A(n137), .B(n185), .C(\send_ppm1/sig_state [2]), 
        .D(\send_ppm1/n91 ), .Q(\send_ppm1/n64 ) );
  OAI212 \send_ppm1/U16  ( .A(\send_ppm1/sig_state [0]), .B(\send_ppm1/n70 ), 
        .C(n130), .Q(\send_ppm1/n66 ) );
  OAI212 \send_ppm1/U13  ( .A(\send_ppm1/n67 ), .B(\send_ppm1/n57 ), .C(
        \send_ppm1/n68 ), .Q(\send_ppm1/n95 ) );
  OAI222 \send_ppm1/U6  ( .A(n129), .B(\send_ppm1/n58 ), .C(n133), .D(
        \send_ppm1/n65 ), .Q(\send_ppm1/n94 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_1  ( .A(
        \send_ppm1/local_counter1/v_val [1]), .B(
        \send_ppm1/local_counter1/v_val [0]), .CO(
        \send_ppm1/local_counter1/add_34/carry [2]), .S(
        \send_ppm1/local_counter1/N7 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_2  ( .A(
        \send_ppm1/local_counter1/v_val [2]), .B(
        \send_ppm1/local_counter1/add_34/carry [2]), .CO(
        \send_ppm1/local_counter1/add_34/carry [3]), .S(
        \send_ppm1/local_counter1/N8 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_3  ( .A(
        \send_ppm1/local_counter1/v_val [3]), .B(
        \send_ppm1/local_counter1/add_34/carry [3]), .CO(
        \send_ppm1/local_counter1/add_34/carry [4]), .S(
        \send_ppm1/local_counter1/N9 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_4  ( .A(
        \send_ppm1/local_counter1/v_val [4]), .B(
        \send_ppm1/local_counter1/add_34/carry [4]), .CO(
        \send_ppm1/local_counter1/add_34/carry [5]), .S(
        \send_ppm1/local_counter1/N10 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_5  ( .A(
        \send_ppm1/local_counter1/v_val [5]), .B(
        \send_ppm1/local_counter1/add_34/carry [5]), .CO(
        \send_ppm1/local_counter1/add_34/carry [6]), .S(
        \send_ppm1/local_counter1/N11 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_6  ( .A(
        \send_ppm1/local_counter1/v_val [6]), .B(
        \send_ppm1/local_counter1/add_34/carry [6]), .CO(
        \send_ppm1/local_counter1/add_34/carry [7]), .S(
        \send_ppm1/local_counter1/N12 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_7  ( .A(
        \send_ppm1/local_counter1/v_val [7]), .B(
        \send_ppm1/local_counter1/add_34/carry [7]), .CO(
        \send_ppm1/local_counter1/add_34/carry [8]), .S(
        \send_ppm1/local_counter1/N13 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_8  ( .A(
        \send_ppm1/local_counter1/v_val [8]), .B(
        \send_ppm1/local_counter1/add_34/carry [8]), .CO(
        \send_ppm1/local_counter1/add_34/carry [9]), .S(
        \send_ppm1/local_counter1/N14 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_9  ( .A(
        \send_ppm1/local_counter1/v_val [9]), .B(
        \send_ppm1/local_counter1/add_34/carry [9]), .CO(
        \send_ppm1/local_counter1/add_34/carry [10]), .S(
        \send_ppm1/local_counter1/N15 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_10  ( .A(
        \send_ppm1/local_counter1/v_val [10]), .B(
        \send_ppm1/local_counter1/add_34/carry [10]), .CO(
        \send_ppm1/local_counter1/add_34/carry [11]), .S(
        \send_ppm1/local_counter1/N16 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_11  ( .A(
        \send_ppm1/local_counter1/v_val [11]), .B(
        \send_ppm1/local_counter1/add_34/carry [11]), .CO(
        \send_ppm1/local_counter1/add_34/carry [12]), .S(
        \send_ppm1/local_counter1/N17 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_12  ( .A(
        \send_ppm1/local_counter1/v_val [12]), .B(
        \send_ppm1/local_counter1/add_34/carry [12]), .CO(
        \send_ppm1/local_counter1/add_34/carry [13]), .S(
        \send_ppm1/local_counter1/N18 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_13  ( .A(
        \send_ppm1/local_counter1/v_val [13]), .B(
        \send_ppm1/local_counter1/add_34/carry [13]), .CO(
        \send_ppm1/local_counter1/add_34/carry [14]), .S(
        \send_ppm1/local_counter1/N19 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_14  ( .A(
        \send_ppm1/local_counter1/v_val [14]), .B(
        \send_ppm1/local_counter1/add_34/carry [14]), .CO(
        \send_ppm1/local_counter1/add_34/carry [15]), .S(
        \send_ppm1/local_counter1/N20 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_15  ( .A(
        \send_ppm1/local_counter1/v_val [15]), .B(
        \send_ppm1/local_counter1/add_34/carry [15]), .CO(
        \send_ppm1/local_counter1/add_34/carry [16]), .S(
        \send_ppm1/local_counter1/N21 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_16  ( .A(
        \send_ppm1/local_counter1/v_val [16]), .B(
        \send_ppm1/local_counter1/add_34/carry [16]), .CO(
        \send_ppm1/local_counter1/add_34/carry [17]), .S(
        \send_ppm1/local_counter1/N22 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_17  ( .A(
        \send_ppm1/local_counter1/v_val [17]), .B(
        \send_ppm1/local_counter1/add_34/carry [17]), .CO(
        \send_ppm1/local_counter1/add_34/carry [18]), .S(
        \send_ppm1/local_counter1/N23 ) );
  ADD22 \send_ppm1/local_counter1/add_34/U1_1_18  ( .A(
        \send_ppm1/local_counter1/v_val [18]), .B(
        \send_ppm1/local_counter1/add_34/carry [18]), .CO(
        \send_ppm1/local_counter1/add_34/carry [19]), .S(
        \send_ppm1/local_counter1/N24 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_2  ( .A(
        \send_ppm1/sig_cyclesTrame2 [2]), .B(\send_ppm1/sig_cyclesTrame3 [2]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [2]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [3]), .S(
        \send_ppm1/dp_cluster_0/N38 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_3  ( .A(
        \send_ppm1/sig_cyclesTrame2 [3]), .B(\send_ppm1/sig_cyclesTrame3 [3]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [3]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [4]), .S(
        \send_ppm1/dp_cluster_0/N39 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_4  ( .A(
        \send_ppm1/sig_cyclesTrame2 [4]), .B(\send_ppm1/sig_cyclesTrame3 [4]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [4]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [5]), .S(
        \send_ppm1/dp_cluster_0/N40 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_5  ( .A(
        \send_ppm1/sig_cyclesTrame2 [5]), .B(\send_ppm1/sig_cyclesTrame3 [5]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [5]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [6]), .S(
        \send_ppm1/dp_cluster_0/N41 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_6  ( .A(
        \send_ppm1/sig_cyclesTrame2 [6]), .B(\send_ppm1/sig_cyclesTrame3 [6]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [6]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [7]), .S(
        \send_ppm1/dp_cluster_0/N42 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_7  ( .A(
        \send_ppm1/sig_cyclesTrame2 [7]), .B(\send_ppm1/sig_cyclesTrame3 [7]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [7]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [8]), .S(
        \send_ppm1/dp_cluster_0/N43 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_8  ( .A(
        \send_ppm1/sig_cyclesTrame2 [8]), .B(\send_ppm1/sig_cyclesTrame3 [8]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [8]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [9]), .S(
        \send_ppm1/dp_cluster_0/N44 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_9  ( .A(
        \send_ppm1/sig_cyclesTrame2 [9]), .B(\send_ppm1/sig_cyclesTrame3 [9]), 
        .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [9]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [10]), .S(
        \send_ppm1/dp_cluster_0/N45 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_10  ( .A(
        \send_ppm1/sig_cyclesTrame2 [10]), .B(\send_ppm1/sig_cyclesTrame3 [10]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [10]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [11]), .S(
        \send_ppm1/dp_cluster_0/N46 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_11  ( .A(
        \send_ppm1/sig_cyclesTrame2 [11]), .B(\send_ppm1/sig_cyclesTrame3 [11]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [11]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [12]), .S(
        \send_ppm1/dp_cluster_0/N47 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_12  ( .A(
        \send_ppm1/sig_cyclesTrame2 [12]), .B(\send_ppm1/sig_cyclesTrame3 [12]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [12]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [13]), .S(
        \send_ppm1/dp_cluster_0/N48 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_13  ( .A(
        \send_ppm1/sig_cyclesTrame2 [13]), .B(\send_ppm1/sig_cyclesTrame3 [13]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [13]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [14]), .S(
        \send_ppm1/dp_cluster_0/N49 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_14  ( .A(
        \send_ppm1/sig_cyclesTrame2 [14]), .B(\send_ppm1/sig_cyclesTrame3 [14]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [14]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [15]), .S(
        \send_ppm1/dp_cluster_0/N50 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/U1_15  ( .A(
        \send_ppm1/sig_cyclesTrame2 [15]), .B(\send_ppm1/sig_cyclesTrame3 [15]), .CI(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [15]), .CO(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [16]), .S(
        \send_ppm1/dp_cluster_0/N51 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_2  ( .A(
        \send_ppm1/dp_cluster_0/N18 ), .B(n201), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [2]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [3]), .S(
        \send_ppm1/dp_cluster_0/N295 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_3  ( .A(
        \send_ppm1/dp_cluster_0/N19 ), .B(n200), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [3]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [4]), .S(
        \send_ppm1/dp_cluster_0/N294 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_4  ( .A(
        \send_ppm1/dp_cluster_0/N20 ), .B(n199), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [4]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [5]), .S(
        \send_ppm1/dp_cluster_0/N293 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_5  ( .A(
        \send_ppm1/dp_cluster_0/N21 ), .B(n198), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [5]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [6]), .S(
        \send_ppm1/dp_cluster_0/N292 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_6  ( .A(
        \send_ppm1/dp_cluster_0/N22 ), .B(n197), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [6]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [7]), .S(
        \send_ppm1/dp_cluster_0/N291 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_7  ( .A(
        \send_ppm1/dp_cluster_0/N23 ), .B(n196), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [7]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [8]), .S(
        \send_ppm1/dp_cluster_0/N290 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_8  ( .A(
        \send_ppm1/dp_cluster_0/N24 ), .B(n195), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [8]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [9]), .S(
        \send_ppm1/dp_cluster_0/N289 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_9  ( .A(
        \send_ppm1/dp_cluster_0/N25 ), .B(n194), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [9]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [10]), .S(
        \send_ppm1/dp_cluster_0/N288 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_10  ( .A(
        \send_ppm1/dp_cluster_0/N26 ), .B(n191), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [10]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [11]), .S(
        \send_ppm1/dp_cluster_0/N287 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_11  ( .A(
        \send_ppm1/dp_cluster_0/N27 ), .B(n190), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [11]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [12]), .S(
        \send_ppm1/dp_cluster_0/N286 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_12  ( .A(
        \send_ppm1/dp_cluster_0/N28 ), .B(n188), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [12]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [13]), .S(
        \send_ppm1/dp_cluster_0/N285 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_13  ( .A(
        \send_ppm1/dp_cluster_0/N29 ), .B(n187), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [13]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [14]), .S(
        \send_ppm1/dp_cluster_0/N284 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_14  ( .A(
        \send_ppm1/dp_cluster_0/N30 ), .B(n186), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [14]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [15]), .S(
        \send_ppm1/dp_cluster_0/N283 ) );
  ADD32 \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/U1_15  ( .A(
        \send_ppm1/dp_cluster_0/N31 ), .B(n47), .CI(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [15]), .CO(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [16]), .S(
        \send_ppm1/dp_cluster_0/N282 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_2  ( .A(
        \send_ppm1/dp_cluster_0/N295 ), .B(n179), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [2]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [3]), .S(
        \send_ppm1/N180 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_3  ( .A(
        \send_ppm1/dp_cluster_0/N294 ), .B(n178), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [3]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [4]), .S(
        \send_ppm1/N181 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_4  ( .A(
        \send_ppm1/dp_cluster_0/N293 ), .B(n177), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [4]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [5]), .S(
        \send_ppm1/N182 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_5  ( .A(
        \send_ppm1/dp_cluster_0/N292 ), .B(n176), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [5]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [6]), .S(
        \send_ppm1/N183 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_6  ( .A(
        \send_ppm1/dp_cluster_0/N291 ), .B(n175), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [6]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [7]), .S(
        \send_ppm1/N184 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_7  ( .A(
        \send_ppm1/dp_cluster_0/N290 ), .B(n174), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [7]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [8]), .S(
        \send_ppm1/N185 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_8  ( .A(
        \send_ppm1/dp_cluster_0/N289 ), .B(n173), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [8]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [9]), .S(
        \send_ppm1/N186 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_9  ( .A(
        \send_ppm1/dp_cluster_0/N288 ), .B(n172), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [9]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [10]), .S(
        \send_ppm1/N187 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_10  ( .A(
        \send_ppm1/dp_cluster_0/N287 ), .B(n169), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [10]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [11]), .S(
        \send_ppm1/N188 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_11  ( .A(
        \send_ppm1/dp_cluster_0/N286 ), .B(n168), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [11]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [12]), .S(
        \send_ppm1/N189 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_12  ( .A(
        \send_ppm1/dp_cluster_0/N285 ), .B(n166), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [12]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [13]), .S(
        \send_ppm1/N190 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_13  ( .A(
        \send_ppm1/dp_cluster_0/N284 ), .B(n165), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [13]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [14]), .S(
        \send_ppm1/N191 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_14  ( .A(
        \send_ppm1/dp_cluster_0/N283 ), .B(n164), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [14]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [15]), .S(
        \send_ppm1/N192 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_15  ( .A(
        \send_ppm1/dp_cluster_0/N282 ), .B(n163), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [15]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [16]), .S(
        \send_ppm1/N193 ) );
  ADD32 \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/U2_16  ( .A(
        \send_ppm1/dp_cluster_0/N281 ), .B(n162), .CI(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [16]), .CO(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [17]), .S(
        \send_ppm1/N194 ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S3_2_5  ( .A(
        \send_ppm1/sig_reg_storage [2]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[1][5] ), .CI(
        \send_ppm1/sig_reg_storage [1]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[2][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[2][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S3_3_5  ( .A(
        \send_ppm1/sig_reg_storage [3]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[2][5] ), .CI(
        \send_ppm1/sig_reg_storage [2]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[3][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[3][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S3_4_5  ( .A(
        \send_ppm1/sig_reg_storage [4]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[3][5] ), .CI(
        \send_ppm1/sig_reg_storage [3]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[4][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S3_5_5  ( .A(
        \send_ppm1/sig_reg_storage [5]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][5] ), .CI(
        \send_ppm1/sig_reg_storage [4]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[5][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S2_5_1  ( .A(
        \send_ppm1/sig_reg_storage [5]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][1] ), .CI(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[1][5] ), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][1] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[5][1] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S3_6_5  ( .A(
        \send_ppm1/sig_reg_storage [6]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][5] ), .CI(
        \send_ppm1/sig_reg_storage [5]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[6][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S2_6_1  ( .A(
        \send_ppm1/sig_reg_storage [6]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[5][1] ), .CI(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[2][5] ), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][1] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[6][1] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S5_5  ( .A(
        \send_ppm1/sig_reg_storage [7]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][5] ), .CI(
        \send_ppm1/sig_reg_storage [6]), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][5] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[7][5] ) );
  ADD32 \send_ppm1/dp_cluster_1/mult_114/S4_1  ( .A(
        \send_ppm1/sig_reg_storage [7]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[6][1] ), .CI(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[3][5] ), .CO(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][1] ), .S(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[7][1] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S3_2_5  ( .A(
        \send_ppm1/sig_reg_storage [10]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[1][5] ), .CI(
        \send_ppm1/sig_reg_storage [9]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[2][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[2][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S3_3_5  ( .A(
        \send_ppm1/sig_reg_storage [11]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[2][5] ), .CI(
        \send_ppm1/sig_reg_storage [10]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[3][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[3][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S3_4_5  ( .A(
        \send_ppm1/sig_reg_storage [12]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[3][5] ), .CI(
        \send_ppm1/sig_reg_storage [11]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[4][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S3_5_5  ( .A(
        \send_ppm1/sig_reg_storage [13]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][5] ), .CI(
        \send_ppm1/sig_reg_storage [12]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[5][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S2_5_1  ( .A(
        \send_ppm1/sig_reg_storage [13]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][1] ), .CI(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[1][5] ), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][1] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[5][1] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S3_6_5  ( .A(
        \send_ppm1/sig_reg_storage [14]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][5] ), .CI(
        \send_ppm1/sig_reg_storage [13]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[6][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S2_6_1  ( .A(
        \send_ppm1/sig_reg_storage [14]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[5][1] ), .CI(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[2][5] ), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][1] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[6][1] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S5_5  ( .A(
        \send_ppm1/sig_reg_storage [15]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][5] ), .CI(
        \send_ppm1/sig_reg_storage [14]), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][5] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[7][5] ) );
  ADD32 \send_ppm1/dp_cluster_2/mult_117/S4_1  ( .A(
        \send_ppm1/sig_reg_storage [15]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[6][1] ), .CI(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[3][5] ), .CO(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][1] ), .S(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[7][1] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S3_2_5  ( .A(
        \send_ppm1/sig_reg_storage [18]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[1][5] ), .CI(
        \send_ppm1/sig_reg_storage [17]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[2][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[2][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S3_3_5  ( .A(
        \send_ppm1/sig_reg_storage [19]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[2][5] ), .CI(
        \send_ppm1/sig_reg_storage [18]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[3][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[3][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S3_4_5  ( .A(
        \send_ppm1/sig_reg_storage [20]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[3][5] ), .CI(
        \send_ppm1/sig_reg_storage [19]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[4][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S3_5_5  ( .A(
        \send_ppm1/sig_reg_storage [21]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][5] ), .CI(
        \send_ppm1/sig_reg_storage [20]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[5][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S2_5_1  ( .A(
        \send_ppm1/sig_reg_storage [21]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][1] ), .CI(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[1][5] ), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][1] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[5][1] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S3_6_5  ( .A(
        \send_ppm1/sig_reg_storage [22]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][5] ), .CI(
        \send_ppm1/sig_reg_storage [21]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[6][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S2_6_1  ( .A(
        \send_ppm1/sig_reg_storage [22]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[5][1] ), .CI(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[2][5] ), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][1] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[6][1] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S5_5  ( .A(
        \send_ppm1/sig_reg_storage [23]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][5] ), .CI(
        \send_ppm1/sig_reg_storage [22]), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][5] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[7][5] ) );
  ADD32 \send_ppm1/dp_cluster_3/mult_120/S4_1  ( .A(
        \send_ppm1/sig_reg_storage [23]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[6][1] ), .CI(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[3][5] ), .CO(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][1] ), .S(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[7][1] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S3_2_5  ( .A(
        \send_ppm1/sig_reg_storage [26]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[1][5] ), .CI(
        \send_ppm1/sig_reg_storage [25]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[2][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[2][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S3_3_5  ( .A(
        \send_ppm1/sig_reg_storage [27]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[2][5] ), .CI(
        \send_ppm1/sig_reg_storage [26]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[3][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[3][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S3_4_5  ( .A(
        \send_ppm1/sig_reg_storage [28]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[3][5] ), .CI(
        \send_ppm1/sig_reg_storage [27]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[4][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S3_5_5  ( .A(
        \send_ppm1/sig_reg_storage [29]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][5] ), .CI(
        \send_ppm1/sig_reg_storage [28]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[5][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S2_5_1  ( .A(
        \send_ppm1/sig_reg_storage [29]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][1] ), .CI(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[1][5] ), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][1] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[5][1] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S3_6_5  ( .A(
        \send_ppm1/sig_reg_storage [30]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][5] ), .CI(
        \send_ppm1/sig_reg_storage [29]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[6][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S2_6_1  ( .A(
        \send_ppm1/sig_reg_storage [30]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[5][1] ), .CI(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[2][5] ), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][1] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[6][1] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S5_5  ( .A(
        \send_ppm1/sig_reg_storage [31]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][5] ), .CI(
        \send_ppm1/sig_reg_storage [30]), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][5] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[7][5] ) );
  ADD32 \send_ppm1/dp_cluster_4/mult_123/S4_1  ( .A(
        \send_ppm1/sig_reg_storage [31]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[6][1] ), .CI(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[3][5] ), .CO(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][1] ), .S(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[7][1] ) );
  DF3 \send_ppm1/sig_state_reg[1]  ( .D(\send_ppm1/n94 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_state [1]), .QN(\send_ppm1/n58 ) );
  DF3 \send_ppm1/current_state_reg[0]  ( .D(\send_ppm1/N81 ), .C(i_clk_top), 
        .Q(\send_ppm1/current_state [0]), .QN(\send_ppm1/n55 ) );
  DF3 \send_ppm1/sig_state_reg[2]  ( .D(\send_ppm1/n95 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_state [2]), .QN(\send_ppm1/n57 ) );
  DF3 \send_ppm1/sig_out_ppm_reg  ( .D(n132), .C(i_clk_top), .Q(o_ppm_top) );
  DF3 \send_ppm1/current_state_reg[2]  ( .D(n131), .C(i_clk_top), .Q(
        \send_ppm1/current_state [2]) );
  DF3 \send_ppm1/current_state_reg[1]  ( .D(\send_ppm1/N82 ), .C(i_clk_top), 
        .Q(\send_ppm1/current_state [1]), .QN(\send_ppm1/n53 ) );
  JK3 \send_ppm1/sig_state_reg[0]  ( .J(\send_ppm1/n69 ), .K(n130), .C(
        i_clk_top), .Q(\send_ppm1/sig_state [0]), .QN(\send_ppm1/n59 ) );
  DF3 \send_ppm1/local_counter1/o_count_reg[0]  ( .D(
        \send_ppm1/local_counter1/N46 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [0]), .QN(n1) );
  DF3 \send_ppm1/local_counter1/o_count_reg[1]  ( .D(
        \send_ppm1/local_counter1/N47 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [1]), .QN(n3) );
  DF3 \send_ppm1/local_counter1/o_count_reg[2]  ( .D(
        \send_ppm1/local_counter1/N48 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [2]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[3]  ( .D(
        \send_ppm1/local_counter1/N49 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [3]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[4]  ( .D(
        \send_ppm1/local_counter1/N50 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [4]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[5]  ( .D(
        \send_ppm1/local_counter1/N51 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [5]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[6]  ( .D(
        \send_ppm1/local_counter1/N52 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [6]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[7]  ( .D(
        \send_ppm1/local_counter1/N53 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [7]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[8]  ( .D(
        \send_ppm1/local_counter1/N54 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [8]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[9]  ( .D(
        \send_ppm1/local_counter1/N55 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [9]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[10]  ( .D(
        \send_ppm1/local_counter1/N56 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [10]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[11]  ( .D(
        \send_ppm1/local_counter1/N57 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [11]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[12]  ( .D(
        \send_ppm1/local_counter1/N58 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [12]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[13]  ( .D(
        \send_ppm1/local_counter1/N59 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [13]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[14]  ( .D(
        \send_ppm1/local_counter1/N60 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [14]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[15]  ( .D(
        \send_ppm1/local_counter1/N61 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [15]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[16]  ( .D(
        \send_ppm1/local_counter1/N62 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [16]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[17]  ( .D(
        \send_ppm1/local_counter1/N63 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [17]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[18]  ( .D(
        \send_ppm1/local_counter1/N64 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [18]) );
  DF3 \send_ppm1/local_counter1/o_count_reg[19]  ( .D(
        \send_ppm1/local_counter1/N65 ), .C(i_clk_top), .Q(
        \send_ppm1/sig_out_local_count [19]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[19]  ( .D(
        \send_ppm1/local_counter1/N65 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [19]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[18]  ( .D(
        \send_ppm1/local_counter1/N64 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [18]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[17]  ( .D(
        \send_ppm1/local_counter1/N63 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [17]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[16]  ( .D(
        \send_ppm1/local_counter1/N62 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [16]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[15]  ( .D(
        \send_ppm1/local_counter1/N61 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [15]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[14]  ( .D(
        \send_ppm1/local_counter1/N60 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [14]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[13]  ( .D(
        \send_ppm1/local_counter1/N59 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [13]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[12]  ( .D(
        \send_ppm1/local_counter1/N58 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [12]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[11]  ( .D(
        \send_ppm1/local_counter1/N57 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [11]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[10]  ( .D(
        \send_ppm1/local_counter1/N56 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [10]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[9]  ( .D(
        \send_ppm1/local_counter1/N55 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [9]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[8]  ( .D(
        \send_ppm1/local_counter1/N54 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [8]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[7]  ( .D(
        \send_ppm1/local_counter1/N53 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [7]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[6]  ( .D(
        \send_ppm1/local_counter1/N52 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [6]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[5]  ( .D(
        \send_ppm1/local_counter1/N51 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [5]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[4]  ( .D(
        \send_ppm1/local_counter1/N50 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [4]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[3]  ( .D(
        \send_ppm1/local_counter1/N49 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [3]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[2]  ( .D(
        \send_ppm1/local_counter1/N48 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [2]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[1]  ( .D(
        \send_ppm1/local_counter1/N47 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [1]) );
  DF3 \send_ppm1/local_counter1/v_val_reg[0]  ( .D(
        \send_ppm1/local_counter1/N46 ), .C(i_clk_top), .Q(
        \send_ppm1/local_counter1/v_val [0]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[6]  ( .D(n123), .E(n127), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [6]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[13]  ( .D(sig_reg[30]), .E(n126), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [13]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[14]  ( .D(sig_reg[30]), .E(n126), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [14]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[22]  ( .D(n123), .E(n125), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [22]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[29]  ( .D(sig_reg[30]), .E(n124), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [29]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[30]  ( .D(sig_reg[30]), .E(n124), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [30]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[5]  ( .D(sig_reg[30]), .E(n127), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [5]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[21]  ( .D(n123), .E(n125), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [21]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[12]  ( .D(sig_reg[30]), .E(n126), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [12]), .QN(n8) );
  DFE1 \send_ppm1/sig_reg_storage_reg[20]  ( .D(sig_reg[30]), .E(n125), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [20]), .QN(n2) );
  DFE1 \send_ppm1/sig_reg_storage_reg[28]  ( .D(n123), .E(n124), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [28]), .QN(n7) );
  DFE1 \send_ppm1/sig_reg_storage_reg[3]  ( .D(n123), .E(n128), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [3]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[10]  ( .D(n123), .E(n127), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [10]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[11]  ( .D(n123), .E(n126), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [11]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[18]  ( .D(sig_reg[30]), .E(n125), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [18]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[19]  ( .D(sig_reg[30]), .E(n125), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [19]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[26]  ( .D(n123), .E(n124), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [26]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[27]  ( .D(sig_reg[30]), .E(n124), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [27]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[4]  ( .D(sig_reg[30]), .E(n127), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [4]), .QN(n4) );
  DFE1 \send_ppm1/sig_reg_storage_reg[2]  ( .D(n123), .E(n128), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [2]) );
  DFE1 \send_ppm1/sig_reg_storage_reg[23]  ( .D(sig_reg[31]), .E(n125), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [23]), .QN(n21) );
  DFE1 \send_ppm1/sig_reg_storage_reg[15]  ( .D(sig_reg[31]), .E(n126), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [15]), .QN(n20) );
  DFE1 \send_ppm1/sig_reg_storage_reg[31]  ( .D(sig_reg[31]), .E(n124), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [31]), .QN(n19) );
  DFE1 \send_ppm1/sig_reg_storage_reg[7]  ( .D(sig_reg[7]), .E(n127), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [7]), .QN(n18) );
  DFE1 \send_ppm1/sig_reg_storage_reg[9]  ( .D(n123), .E(n127), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [9]), .QN(n17) );
  DFE1 \send_ppm1/sig_reg_storage_reg[17]  ( .D(n123), .E(n126), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [17]), .QN(n16) );
  DFE1 \send_ppm1/sig_reg_storage_reg[25]  ( .D(n123), .E(n124), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [25]), .QN(n15) );
  DFE1 \send_ppm1/sig_reg_storage_reg[8]  ( .D(sig_reg[30]), .E(n127), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [8]), .QN(n14) );
  DFE1 \send_ppm1/sig_reg_storage_reg[16]  ( .D(sig_reg[30]), .E(n126), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [16]), .QN(n13) );
  DFE1 \send_ppm1/sig_reg_storage_reg[1]  ( .D(sig_reg[30]), .E(n128), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [1]), .QN(n6) );
  DFE1 \send_ppm1/sig_reg_storage_reg[24]  ( .D(sig_reg[30]), .E(n125), .C(
        i_clk_top), .Q(\send_ppm1/sig_reg_storage [24]), .QN(n22) );
  DFE1 \send_ppm1/sig_reg_storage_reg[0]  ( .D(n123), .E(n128), .C(i_clk_top), 
        .Q(\send_ppm1/sig_reg_storage [0]), .QN(n9) );
  NOR21 U1 ( .A(n121), .B(n24), .Q(\send_ppm1/local_counter1/N65 ) );
  MUX22 U2 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[5][5] ), .B(n150), .S(
        \send_ppm1/dp_cluster_1/mult_114/A2[8] ), .Q(n5) );
  MUX22 U3 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[5][5] ), .B(n192), .S(
        \send_ppm1/dp_cluster_4/mult_123/A2[8] ), .Q(n10) );
  MUX22 U4 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[5][5] ), .B(n182), .S(
        \send_ppm1/dp_cluster_3/mult_120/A2[8] ), .Q(n11) );
  MUX22 U5 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[5][5] ), .B(n170), .S(
        \send_ppm1/dp_cluster_2/mult_117/A2[8] ), .Q(n12) );
  XNR21 U6 ( .A(n143), .B(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [18]), .Q(
        \send_ppm1/dp_cluster_0/N279 ) );
  XNR21 U7 ( .A(\send_ppm1/dp_cluster_0/N279 ), .B(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [18]), .Q(
        \send_ppm1/N196 ) );
  INV3 U8 ( .A(\send_ppm1/dp_cluster_0/N48 ), .Q(n166) );
  NOR21 U9 ( .A(\send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [18]), .B(
        \send_ppm1/dp_cluster_0/N279 ), .Q(n55) );
  NOR21 U10 ( .A(\send_ppm1/sig_cyclesTrame1 [12]), .B(n60), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [13]) );
  INV3 U11 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [12]), .Q(
        n60) );
  INV3 U12 ( .A(n53), .Q(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [19]) );
  NOR21 U13 ( .A(\send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [18]), 
        .B(n143), .Q(n53) );
  XNR21 U14 ( .A(n143), .B(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [17]), .Q(
        \send_ppm1/dp_cluster_0/N280 ) );
  INV3 U15 ( .A(\send_ppm1/sig_cyclesTrame4 [12]), .Q(n188) );
  XOR21 U16 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [12]), 
        .B(n146), .Q(\send_ppm1/dp_cluster_0/N28 ) );
  INV3 U17 ( .A(\send_ppm1/dp_cluster_0/N45 ), .Q(n172) );
  INV3 U18 ( .A(\send_ppm1/dp_cluster_0/N46 ), .Q(n169) );
  INV3 U19 ( .A(\send_ppm1/dp_cluster_0/N47 ), .Q(n168) );
  INV3 U20 ( .A(\send_ppm1/dp_cluster_0/N49 ), .Q(n165) );
  INV3 U21 ( .A(n54), .Q(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [18]) );
  NOR21 U22 ( .A(\send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [17]), 
        .B(\send_ppm1/dp_cluster_0/N280 ), .Q(n54) );
  INV3 U23 ( .A(n52), .Q(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [18]) );
  NOR21 U24 ( .A(\send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [17]), 
        .B(n143), .Q(n52) );
  NOR21 U25 ( .A(\send_ppm1/sig_cyclesTrame1 [13]), .B(n61), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [14]) );
  INV3 U26 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [13]), .Q(
        n61) );
  NOR21 U27 ( .A(\send_ppm1/sig_cyclesTrame1 [11]), .B(n59), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [12]) );
  INV3 U28 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [11]), .Q(
        n59) );
  NOR21 U29 ( .A(\send_ppm1/sig_cyclesTrame1 [10]), .B(n27), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [11]) );
  INV3 U30 ( .A(\send_ppm1/sig_cyclesTrame1 [12]), .Q(n146) );
  INV3 U31 ( .A(n27), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [10]) );
  NOR21 U32 ( .A(n152), .B(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [9]), .Q(n27) );
  INV3 U33 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [16]), .Q(
        n143) );
  INV3 U34 ( .A(\send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [16]), .Q(
        n162) );
  XNR21 U35 ( .A(n143), .B(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [16]), .Q(
        \send_ppm1/dp_cluster_0/N281 ) );
  INV3 U36 ( .A(\send_ppm1/sig_cyclesTrame4 [10]), .Q(n191) );
  XOR21 U37 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [10]), 
        .B(n149), .Q(\send_ppm1/dp_cluster_0/N26 ) );
  INV3 U38 ( .A(\send_ppm1/sig_cyclesTrame4 [9]), .Q(n194) );
  XNR21 U39 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [9]), .B(
        n152), .Q(\send_ppm1/dp_cluster_0/N25 ) );
  INV3 U40 ( .A(\send_ppm1/sig_cyclesTrame4 [13]), .Q(n187) );
  XOR21 U41 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [13]), 
        .B(n145), .Q(\send_ppm1/dp_cluster_0/N29 ) );
  INV3 U42 ( .A(\send_ppm1/sig_cyclesTrame4 [11]), .Q(n190) );
  XOR21 U43 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [11]), 
        .B(n148), .Q(\send_ppm1/dp_cluster_0/N27 ) );
  INV3 U44 ( .A(\send_ppm1/dp_cluster_0/N41 ), .Q(n176) );
  INV3 U45 ( .A(\send_ppm1/dp_cluster_0/N42 ), .Q(n175) );
  INV3 U46 ( .A(\send_ppm1/dp_cluster_0/N43 ), .Q(n174) );
  INV3 U47 ( .A(\send_ppm1/dp_cluster_0/N44 ), .Q(n173) );
  INV3 U48 ( .A(\send_ppm1/dp_cluster_0/N50 ), .Q(n164) );
  INV3 U49 ( .A(\send_ppm1/dp_cluster_0/N51 ), .Q(n163) );
  INV3 U50 ( .A(n51), .Q(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [17]) );
  NOR21 U51 ( .A(\send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [16]), 
        .B(n143), .Q(n51) );
  XOR21 U52 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [12]), .B(
        \send_ppm1/dp_cluster_2/N250 ), .Q(\send_ppm1/sig_cyclesTrame2 [12])
         );
  XOR21 U53 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [12]), .B(
        \send_ppm1/dp_cluster_3/N235 ), .Q(\send_ppm1/sig_cyclesTrame3 [12])
         );
  XOR21 U54 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [12]), .B(
        \send_ppm1/dp_cluster_1/N265 ), .Q(\send_ppm1/sig_cyclesTrame1 [12])
         );
  XOR21 U55 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [12]), .B(
        \send_ppm1/dp_cluster_4/N220 ), .Q(\send_ppm1/sig_cyclesTrame4 [12])
         );
  NOR21 U56 ( .A(\send_ppm1/sig_cyclesTrame1 [5]), .B(n58), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [6]) );
  INV3 U57 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [5]), .Q(
        n58) );
  NOR21 U58 ( .A(\send_ppm1/sig_cyclesTrame1 [8]), .B(n26), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [9]) );
  NOR21 U59 ( .A(n102), .B(n103), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [13]) );
  INV3 U60 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [12]), .Q(n102) );
  INV3 U61 ( .A(\send_ppm1/dp_cluster_3/N235 ), .Q(n103) );
  NOR21 U62 ( .A(\send_ppm1/sig_cyclesTrame1 [14]), .B(n62), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [15]) );
  INV3 U63 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [14]), .Q(
        n62) );
  INV3 U64 ( .A(\send_ppm1/sig_cyclesTrame1 [9]), .Q(n152) );
  INV3 U65 ( .A(\send_ppm1/sig_cyclesTrame1 [13]), .Q(n145) );
  INV3 U66 ( .A(\send_ppm1/sig_cyclesTrame1 [11]), .Q(n148) );
  INV3 U67 ( .A(\send_ppm1/sig_cyclesTrame1 [10]), .Q(n149) );
  NOR21 U68 ( .A(n74), .B(n75), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [13]) );
  INV3 U69 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [12]), .Q(n74) );
  INV3 U70 ( .A(\send_ppm1/dp_cluster_1/N265 ), .Q(n75) );
  INV3 U71 ( .A(n25), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [7]) );
  NOR21 U72 ( .A(n155), .B(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [6]), .Q(n25) );
  INV3 U73 ( .A(n26), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [8]) );
  NOR21 U74 ( .A(n154), .B(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [7]), .Q(n26) );
  NOR21 U75 ( .A(n88), .B(n89), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [13]) );
  INV3 U76 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [12]), .Q(n88) );
  INV3 U77 ( .A(\send_ppm1/dp_cluster_2/N250 ), .Q(n89) );
  NOR21 U78 ( .A(n116), .B(n117), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [13]) );
  INV3 U79 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [12]), .Q(n116) );
  INV3 U80 ( .A(\send_ppm1/dp_cluster_4/N220 ), .Q(n117) );
  NOR21 U81 ( .A(\send_ppm1/sig_cyclesTrame1 [15]), .B(n63), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [16]) );
  INV3 U82 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [15]), .Q(
        n63) );
  XOR21 U83 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [15]), 
        .B(n32), .Q(\send_ppm1/dp_cluster_0/N31 ) );
  INV3 U84 ( .A(\send_ppm1/sig_cyclesTrame4 [6]), .Q(n197) );
  XNR21 U85 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [6]), .B(
        n155), .Q(\send_ppm1/dp_cluster_0/N22 ) );
  INV3 U86 ( .A(\send_ppm1/sig_cyclesTrame4 [14]), .Q(n186) );
  XOR21 U87 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [14]), 
        .B(n144), .Q(\send_ppm1/dp_cluster_0/N30 ) );
  INV3 U88 ( .A(\send_ppm1/sig_cyclesTrame4 [5]), .Q(n198) );
  XOR21 U89 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [5]), .B(
        n156), .Q(\send_ppm1/dp_cluster_0/N21 ) );
  INV3 U90 ( .A(\send_ppm1/sig_cyclesTrame4 [7]), .Q(n196) );
  XNR21 U91 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [7]), .B(
        n154), .Q(\send_ppm1/dp_cluster_0/N23 ) );
  INV3 U92 ( .A(\send_ppm1/sig_cyclesTrame4 [8]), .Q(n195) );
  XOR21 U93 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [8]), .B(
        n153), .Q(\send_ppm1/dp_cluster_0/N24 ) );
  INV3 U94 ( .A(\send_ppm1/dp_cluster_0/N39 ), .Q(n178) );
  INV3 U95 ( .A(\send_ppm1/dp_cluster_0/N40 ), .Q(n177) );
  INV3 U96 ( .A(\send_ppm1/N198 ), .Q(n141) );
  XOR21 U97 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [11]), .B(
        \send_ppm1/dp_cluster_2/N251 ), .Q(\send_ppm1/sig_cyclesTrame2 [11])
         );
  XOR21 U98 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [13]), .B(
        \send_ppm1/dp_cluster_3/N234 ), .Q(\send_ppm1/sig_cyclesTrame3 [13])
         );
  XOR21 U99 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [11]), .B(
        \send_ppm1/dp_cluster_3/N236 ), .Q(\send_ppm1/sig_cyclesTrame3 [11])
         );
  XOR21 U100 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [9]), .B(
        \send_ppm1/dp_cluster_1/N268 ), .Q(\send_ppm1/sig_cyclesTrame1 [9]) );
  XOR21 U101 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [13]), .B(
        \send_ppm1/dp_cluster_1/N264 ), .Q(\send_ppm1/sig_cyclesTrame1 [13])
         );
  XOR21 U102 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [11]), .B(
        \send_ppm1/dp_cluster_1/N266 ), .Q(\send_ppm1/sig_cyclesTrame1 [11])
         );
  XOR21 U103 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [11]), .B(
        \send_ppm1/dp_cluster_4/N221 ), .Q(\send_ppm1/sig_cyclesTrame4 [11])
         );
  XOR21 U104 ( .A(n246), .B(n147), .Q(\send_ppm1/dp_cluster_1/N265 ) );
  XOR21 U105 ( .A(n228), .B(n189), .Q(\send_ppm1/dp_cluster_4/N220 ) );
  XOR21 U106 ( .A(n234), .B(n181), .Q(\send_ppm1/dp_cluster_3/N235 ) );
  XOR21 U107 ( .A(n240), .B(n167), .Q(\send_ppm1/dp_cluster_2/N250 ) );
  XNR21 U108 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [10]), .B(n5), .Q(
        \send_ppm1/sig_cyclesTrame1 [10]) );
  NOR21 U109 ( .A(n76), .B(n77), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [14]) );
  INV3 U110 ( .A(\send_ppm1/dp_cluster_1/N264 ), .Q(n77) );
  INV3 U111 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [13]), .Q(n76) );
  NOR21 U112 ( .A(n46), .B(n115), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [12]) );
  INV3 U113 ( .A(\send_ppm1/dp_cluster_4/N221 ), .Q(n115) );
  NOR21 U114 ( .A(n41), .B(n101), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [12]) );
  INV3 U115 ( .A(\send_ppm1/dp_cluster_3/N236 ), .Q(n101) );
  NOR21 U116 ( .A(n36), .B(n87), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [12]) );
  INV3 U117 ( .A(\send_ppm1/dp_cluster_2/N251 ), .Q(n87) );
  NOR21 U118 ( .A(\send_ppm1/sig_cyclesTrame1 [4]), .B(n57), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [5]) );
  INV3 U119 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [4]), .Q(
        n57) );
  INV3 U120 ( .A(\send_ppm1/sig_cyclesTrame1 [7]), .Q(n154) );
  INV3 U121 ( .A(\send_ppm1/sig_cyclesTrame1 [8]), .Q(n153) );
  INV3 U122 ( .A(\send_ppm1/sig_cyclesTrame1 [5]), .Q(n156) );
  INV3 U123 ( .A(\send_ppm1/sig_cyclesTrame1 [6]), .Q(n155) );
  INV3 U124 ( .A(\send_ppm1/sig_cyclesTrame1 [14]), .Q(n144) );
  NOR21 U125 ( .A(n71), .B(n72), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [10]) );
  INV3 U126 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [9]), .Q(n71) );
  INV3 U127 ( .A(\send_ppm1/dp_cluster_1/N268 ), .Q(n72) );
  NOR21 U128 ( .A(n31), .B(n73), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [12]) );
  INV3 U129 ( .A(\send_ppm1/dp_cluster_1/N266 ), .Q(n73) );
  INV3 U130 ( .A(n31), .Q(\send_ppm1/dp_cluster_1/sub_114_cf/carry [11]) );
  NOR21 U131 ( .A(n5), .B(\send_ppm1/dp_cluster_1/sub_114_cf/carry [10]), .Q(
        n31) );
  XOR21 U132 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [13]), .B(
        \send_ppm1/dp_cluster_2/N249 ), .Q(\send_ppm1/sig_cyclesTrame2 [13])
         );
  XOR21 U133 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [9]), .B(
        \send_ppm1/dp_cluster_2/N253 ), .Q(\send_ppm1/sig_cyclesTrame2 [9]) );
  XOR21 U134 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [9]), .B(
        \send_ppm1/dp_cluster_3/N238 ), .Q(\send_ppm1/sig_cyclesTrame3 [9]) );
  XNR21 U135 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [10]), .B(n12), .Q(
        \send_ppm1/sig_cyclesTrame2 [10]) );
  XNR21 U136 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [10]), .B(n11), .Q(
        \send_ppm1/sig_cyclesTrame3 [10]) );
  XOR21 U137 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [13]), .B(
        \send_ppm1/dp_cluster_4/N219 ), .Q(\send_ppm1/sig_cyclesTrame4 [13])
         );
  XOR21 U138 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [9]), .B(
        \send_ppm1/dp_cluster_4/N223 ), .Q(\send_ppm1/sig_cyclesTrame4 [9]) );
  XNR21 U139 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [10]), .B(n10), .Q(
        \send_ppm1/sig_cyclesTrame4 [10]) );
  NOR21 U140 ( .A(n99), .B(n100), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [10]) );
  INV3 U141 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [9]), .Q(n99) );
  INV3 U142 ( .A(\send_ppm1/dp_cluster_3/N238 ), .Q(n100) );
  NOR21 U143 ( .A(n85), .B(n86), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [10]) );
  INV3 U144 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [9]), .Q(n85) );
  INV3 U145 ( .A(\send_ppm1/dp_cluster_2/N253 ), .Q(n86) );
  NOR21 U146 ( .A(n118), .B(n119), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [14]) );
  INV3 U147 ( .A(\send_ppm1/dp_cluster_4/N219 ), .Q(n119) );
  INV3 U148 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [13]), .Q(n118) );
  NOR21 U149 ( .A(n104), .B(n105), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [14]) );
  INV3 U150 ( .A(\send_ppm1/dp_cluster_3/N234 ), .Q(n105) );
  INV3 U151 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [13]), .Q(n104) );
  NOR21 U152 ( .A(n90), .B(n91), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [14]) );
  INV3 U153 ( .A(\send_ppm1/dp_cluster_2/N249 ), .Q(n91) );
  INV3 U154 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [13]), .Q(n90) );
  INV3 U155 ( .A(n46), .Q(\send_ppm1/dp_cluster_4/sub_123_cf/carry [11]) );
  NOR21 U156 ( .A(n10), .B(\send_ppm1/dp_cluster_4/sub_123_cf/carry [10]), .Q(
        n46) );
  INV3 U157 ( .A(n41), .Q(\send_ppm1/dp_cluster_3/sub_120_cf/carry [11]) );
  NOR21 U158 ( .A(n11), .B(\send_ppm1/dp_cluster_3/sub_120_cf/carry [10]), .Q(
        n41) );
  INV3 U159 ( .A(n36), .Q(\send_ppm1/dp_cluster_2/sub_117_cf/carry [11]) );
  NOR21 U160 ( .A(n12), .B(\send_ppm1/dp_cluster_2/sub_117_cf/carry [10]), .Q(
        n36) );
  NOR21 U161 ( .A(n113), .B(n114), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [10]) );
  INV3 U162 ( .A(\send_ppm1/dp_cluster_4/N223 ), .Q(n114) );
  INV3 U163 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [9]), .Q(n113) );
  BUF2 U164 ( .A(n138), .Q(n124) );
  BUF2 U165 ( .A(n138), .Q(n125) );
  BUF2 U166 ( .A(n138), .Q(n126) );
  BUF2 U167 ( .A(n138), .Q(n127) );
  BUF2 U168 ( .A(n138), .Q(n128) );
  NOR40 U169 ( .A(n142), .B(n275), .C(n274), .D(n273), .Q(\send_ppm1/N198 ) );
  NAND31 U170 ( .A(n270), .B(n269), .C(n268), .Q(n274) );
  NAND22 U171 ( .A(n272), .B(n271), .Q(n273) );
  INV3 U172 ( .A(n261), .Q(n142) );
  NAND41 U173 ( .A(n161), .B(n267), .C(n266), .D(n265), .Q(n275) );
  NAND22 U174 ( .A(n3), .B(\send_ppm1/N179 ), .Q(n267) );
  INV3 U175 ( .A(n262), .Q(n161) );
  NOR21 U176 ( .A(n264), .B(n263), .Q(n265) );
  NOR40 U177 ( .A(n260), .B(n259), .C(n258), .D(n257), .Q(n261) );
  NAND31 U178 ( .A(n249), .B(n248), .C(n247), .Q(n260) );
  NAND22 U179 ( .A(n251), .B(n250), .Q(n259) );
  NAND31 U180 ( .A(n254), .B(n253), .C(n252), .Q(n258) );
  NOR21 U181 ( .A(\send_ppm1/sig_cyclesTrame1 [3]), .B(n56), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [4]) );
  INV3 U182 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [3]), .Q(
        n56) );
  INV3 U183 ( .A(\send_ppm1/sig_cyclesTrame4 [3]), .Q(n200) );
  XOR21 U184 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [3]), 
        .B(n158), .Q(\send_ppm1/dp_cluster_0/N19 ) );
  INV3 U185 ( .A(\send_ppm1/sig_cyclesTrame4 [4]), .Q(n199) );
  XOR21 U186 ( .A(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [4]), 
        .B(n157), .Q(\send_ppm1/dp_cluster_0/N20 ) );
  INV3 U187 ( .A(n50), .Q(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [2]) );
  INV3 U188 ( .A(\send_ppm1/dp_cluster_0/N38 ), .Q(n179) );
  NOR21 U189 ( .A(n23), .B(\send_ppm1/dp_cluster_0/N296 ), .Q(n50) );
  BUF2 U190 ( .A(\send_ppm1/local_counter1/n22 ), .Q(n121) );
  BUF2 U191 ( .A(\send_ppm1/local_counter1/n22 ), .Q(n120) );
  INV3 U192 ( .A(\send_ppm1/sig_cyclesTrame1 [2]), .Q(n159) );
  INV3 U193 ( .A(\send_ppm1/sig_cyclesTrame1 [3]), .Q(n158) );
  INV3 U194 ( .A(\send_ppm1/sig_cyclesTrame1 [4]), .Q(n157) );
  NOR21 U195 ( .A(n121), .B(n206), .Q(\send_ppm1/local_counter1/N63 ) );
  INV3 U196 ( .A(\send_ppm1/local_counter1/N23 ), .Q(n206) );
  NOR21 U197 ( .A(n121), .B(n208), .Q(\send_ppm1/local_counter1/N61 ) );
  INV3 U198 ( .A(\send_ppm1/local_counter1/N21 ), .Q(n208) );
  NOR21 U199 ( .A(n121), .B(n210), .Q(\send_ppm1/local_counter1/N59 ) );
  INV3 U200 ( .A(\send_ppm1/local_counter1/N19 ), .Q(n210) );
  NOR21 U201 ( .A(n121), .B(n212), .Q(\send_ppm1/local_counter1/N57 ) );
  INV3 U202 ( .A(\send_ppm1/local_counter1/N17 ), .Q(n212) );
  NOR21 U203 ( .A(n121), .B(n214), .Q(\send_ppm1/local_counter1/N55 ) );
  INV3 U204 ( .A(\send_ppm1/local_counter1/N15 ), .Q(n214) );
  NOR21 U205 ( .A(n121), .B(n216), .Q(\send_ppm1/local_counter1/N53 ) );
  INV3 U206 ( .A(\send_ppm1/local_counter1/N13 ), .Q(n216) );
  NOR21 U207 ( .A(n120), .B(n217), .Q(\send_ppm1/local_counter1/N52 ) );
  INV3 U208 ( .A(\send_ppm1/local_counter1/N12 ), .Q(n217) );
  NOR21 U209 ( .A(n120), .B(n218), .Q(\send_ppm1/local_counter1/N51 ) );
  INV3 U210 ( .A(\send_ppm1/local_counter1/N11 ), .Q(n218) );
  NOR21 U211 ( .A(n120), .B(n219), .Q(\send_ppm1/local_counter1/N50 ) );
  INV3 U212 ( .A(\send_ppm1/local_counter1/N10 ), .Q(n219) );
  NOR21 U213 ( .A(n120), .B(n220), .Q(\send_ppm1/local_counter1/N49 ) );
  INV3 U214 ( .A(\send_ppm1/local_counter1/N9 ), .Q(n220) );
  NOR21 U215 ( .A(n120), .B(n221), .Q(\send_ppm1/local_counter1/N48 ) );
  INV3 U216 ( .A(\send_ppm1/local_counter1/N8 ), .Q(n221) );
  NOR21 U217 ( .A(n120), .B(n222), .Q(\send_ppm1/local_counter1/N47 ) );
  INV3 U218 ( .A(\send_ppm1/local_counter1/N7 ), .Q(n222) );
  XOR21 U219 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [5]), .B(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[4][1] ), .Q(
        \send_ppm1/sig_cyclesTrame2 [5]) );
  XOR21 U220 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [8]), .B(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[7][1] ), .Q(
        \send_ppm1/sig_cyclesTrame3 [8]) );
  XOR21 U221 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [5]), .B(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[4][1] ), .Q(
        \send_ppm1/sig_cyclesTrame3 [5]) );
  XOR21 U222 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [8]), .B(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[7][1] ), .Q(
        \send_ppm1/sig_cyclesTrame1 [8]) );
  XOR21 U223 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [8]), .B(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[7][1] ), .Q(
        \send_ppm1/sig_cyclesTrame4 [8]) );
  XOR21 U224 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [5]), .B(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[4][1] ), .Q(
        \send_ppm1/sig_cyclesTrame1 [5]) );
  XOR21 U225 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [5]), .B(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[4][1] ), .Q(
        \send_ppm1/sig_cyclesTrame4 [5]) );
  XOR21 U226 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [7]), .B(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[6][1] ), .Q(
        \send_ppm1/sig_cyclesTrame1 [7]) );
  XOR21 U227 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [7]), .B(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[6][1] ), .Q(
        \send_ppm1/sig_cyclesTrame4 [7]) );
  XOR21 U228 ( .A(\send_ppm1/dp_cluster_1/mult_114/A1[11] ), .B(n245), .Q(
        \send_ppm1/dp_cluster_1/N264 ) );
  NOR21 U229 ( .A(n147), .B(n246), .Q(n245) );
  XOR21 U230 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[4][5] ), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][1] ), .Q(
        \send_ppm1/dp_cluster_1/N268 ) );
  XNR21 U231 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [14]), .B(
        \send_ppm1/dp_cluster_1/N263 ), .Q(\send_ppm1/sig_cyclesTrame1 [14])
         );
  XNR21 U232 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [6]), .B(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[5][1] ), .Q(
        \send_ppm1/sig_cyclesTrame1 [6]) );
  XNR21 U233 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [6]), .B(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[5][1] ), .Q(
        \send_ppm1/sig_cyclesTrame4 [6]) );
  XOR21 U234 ( .A(n151), .B(\send_ppm1/dp_cluster_1/mult_114/SUMB[6][5] ), .Q(
        \send_ppm1/dp_cluster_1/N266 ) );
  XOR21 U235 ( .A(n193), .B(\send_ppm1/dp_cluster_4/mult_123/SUMB[6][5] ), .Q(
        \send_ppm1/dp_cluster_4/N221 ) );
  XOR21 U236 ( .A(n183), .B(\send_ppm1/dp_cluster_3/mult_120/SUMB[6][5] ), .Q(
        \send_ppm1/dp_cluster_3/N236 ) );
  XOR21 U237 ( .A(n171), .B(\send_ppm1/dp_cluster_2/mult_117/SUMB[6][5] ), .Q(
        \send_ppm1/dp_cluster_2/N251 ) );
  NAND22 U238 ( .A(n151), .B(\send_ppm1/dp_cluster_1/mult_114/SUMB[6][5] ), 
        .Q(n246) );
  NOR21 U239 ( .A(n29), .B(n67), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [6]) );
  INV3 U240 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[4][1] ), .Q(n67) );
  NOR21 U241 ( .A(n64), .B(n65), .Q(\send_ppm1/dp_cluster_1/mult_114/A2[8] )
         );
  INV3 U242 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[4][5] ), .Q(n65) );
  INV3 U243 ( .A(\send_ppm1/dp_cluster_1/mult_114/CARRYB[7][1] ), .Q(n64) );
  NOR21 U244 ( .A(n69), .B(n70), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [9]) );
  INV3 U245 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [8]), .Q(n69) );
  INV3 U246 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[7][1] ), .Q(n70) );
  NOR21 U247 ( .A(n30), .B(n68), .Q(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [8]) );
  INV3 U248 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[6][1] ), .Q(n68) );
  INV3 U249 ( .A(n49), .Q(
        \send_ppm1/dp_cluster_0/add_3_root_sub_235_cf/carry [2]) );
  NOR21 U250 ( .A(n13), .B(n14), .Q(n49) );
  INV3 U251 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[7][5] ), .Q(n147) );
  INV3 U252 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[7][5] ), .Q(n189) );
  INV3 U253 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[7][5] ), .Q(n181) );
  INV3 U254 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[7][5] ), .Q(n167) );
  INV3 U255 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[5][5] ), .Q(n150) );
  INV3 U256 ( .A(n241), .Q(n151) );
  NAND22 U257 ( .A(\send_ppm1/dp_cluster_1/mult_114/A2[8] ), .B(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[5][5] ), .Q(n241) );
  BUF2 U258 ( .A(\send_ppm1/local_counter1/n22 ), .Q(n122) );
  XOR21 U259 ( .A(n14), .B(n13), .Q(n23) );
  INV3 U260 ( .A(n30), .Q(\send_ppm1/dp_cluster_1/sub_114_cf/carry [7]) );
  NOR21 U261 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[5][1] ), .B(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [6]), .Q(n30) );
  NOR21 U262 ( .A(n122), .B(n205), .Q(\send_ppm1/local_counter1/N64 ) );
  INV3 U263 ( .A(\send_ppm1/local_counter1/N24 ), .Q(n205) );
  NOR21 U264 ( .A(n122), .B(n207), .Q(\send_ppm1/local_counter1/N62 ) );
  INV3 U265 ( .A(\send_ppm1/local_counter1/N22 ), .Q(n207) );
  NOR21 U266 ( .A(n122), .B(n209), .Q(\send_ppm1/local_counter1/N60 ) );
  INV3 U267 ( .A(\send_ppm1/local_counter1/N20 ), .Q(n209) );
  NOR21 U268 ( .A(n122), .B(n211), .Q(\send_ppm1/local_counter1/N58 ) );
  INV3 U269 ( .A(\send_ppm1/local_counter1/N18 ), .Q(n211) );
  NOR21 U270 ( .A(n122), .B(n213), .Q(\send_ppm1/local_counter1/N56 ) );
  INV3 U271 ( .A(\send_ppm1/local_counter1/N16 ), .Q(n213) );
  NOR21 U272 ( .A(n122), .B(n215), .Q(\send_ppm1/local_counter1/N54 ) );
  INV3 U273 ( .A(\send_ppm1/local_counter1/N14 ), .Q(n215) );
  XOR21 U274 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [8]), .B(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[7][1] ), .Q(
        \send_ppm1/sig_cyclesTrame2 [8]) );
  XOR21 U275 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [7]), .B(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[6][1] ), .Q(
        \send_ppm1/sig_cyclesTrame2 [7]) );
  XOR21 U276 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [7]), .B(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[6][1] ), .Q(
        \send_ppm1/sig_cyclesTrame3 [7]) );
  XNR21 U277 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [14]), .B(
        \send_ppm1/dp_cluster_2/N248 ), .Q(\send_ppm1/sig_cyclesTrame2 [14])
         );
  XNR21 U278 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [6]), .B(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[5][1] ), .Q(
        \send_ppm1/sig_cyclesTrame2 [6]) );
  XNR21 U279 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [14]), .B(
        \send_ppm1/dp_cluster_3/N233 ), .Q(\send_ppm1/sig_cyclesTrame3 [14])
         );
  XNR21 U280 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [6]), .B(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[5][1] ), .Q(
        \send_ppm1/sig_cyclesTrame3 [6]) );
  XOR21 U281 ( .A(\send_ppm1/dp_cluster_4/mult_123/A1[11] ), .B(n227), .Q(
        \send_ppm1/dp_cluster_4/N219 ) );
  NOR21 U282 ( .A(n189), .B(n228), .Q(n227) );
  XOR21 U283 ( .A(\send_ppm1/dp_cluster_3/mult_120/A1[11] ), .B(n233), .Q(
        \send_ppm1/dp_cluster_3/N234 ) );
  NOR21 U284 ( .A(n181), .B(n234), .Q(n233) );
  XOR21 U285 ( .A(\send_ppm1/dp_cluster_2/mult_117/A1[11] ), .B(n239), .Q(
        \send_ppm1/dp_cluster_2/N249 ) );
  NOR21 U286 ( .A(n167), .B(n240), .Q(n239) );
  XOR21 U287 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[4][5] ), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][1] ), .Q(
        \send_ppm1/dp_cluster_4/N223 ) );
  XOR21 U288 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[4][5] ), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][1] ), .Q(
        \send_ppm1/dp_cluster_3/N238 ) );
  XOR21 U289 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[4][5] ), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][1] ), .Q(
        \send_ppm1/dp_cluster_2/N253 ) );
  XNR21 U290 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [14]), .B(
        \send_ppm1/dp_cluster_4/N218 ), .Q(\send_ppm1/sig_cyclesTrame4 [14])
         );
  NAND22 U291 ( .A(n193), .B(\send_ppm1/dp_cluster_4/mult_123/SUMB[6][5] ), 
        .Q(n228) );
  NAND22 U292 ( .A(n183), .B(\send_ppm1/dp_cluster_3/mult_120/SUMB[6][5] ), 
        .Q(n234) );
  NAND22 U293 ( .A(n171), .B(\send_ppm1/dp_cluster_2/mult_117/SUMB[6][5] ), 
        .Q(n240) );
  NOR21 U294 ( .A(n44), .B(n109), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [6]) );
  INV3 U295 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[4][1] ), .Q(n109) );
  NOR21 U296 ( .A(n39), .B(n95), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [6]) );
  INV3 U297 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[4][1] ), .Q(n95) );
  NOR21 U298 ( .A(n34), .B(n81), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [6]) );
  INV3 U299 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[4][1] ), .Q(n81) );
  NOR21 U300 ( .A(n106), .B(n107), .Q(\send_ppm1/dp_cluster_4/mult_123/A2[8] )
         );
  INV3 U301 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[4][5] ), .Q(n107) );
  INV3 U302 ( .A(\send_ppm1/dp_cluster_4/mult_123/CARRYB[7][1] ), .Q(n106) );
  NOR21 U303 ( .A(n111), .B(n112), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [9]) );
  INV3 U304 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [8]), .Q(n111) );
  INV3 U305 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[7][1] ), .Q(n112) );
  NOR21 U306 ( .A(n97), .B(n98), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [9]) );
  INV3 U307 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [8]), .Q(n97) );
  INV3 U308 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[7][1] ), .Q(n98) );
  NOR21 U309 ( .A(n83), .B(n84), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [9]) );
  INV3 U310 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [8]), .Q(n83) );
  INV3 U311 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[7][1] ), .Q(n84) );
  NOR21 U312 ( .A(n45), .B(n110), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [8]) );
  INV3 U313 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[6][1] ), .Q(n110) );
  NOR21 U314 ( .A(n40), .B(n96), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [8]) );
  INV3 U315 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[6][1] ), .Q(n96) );
  NOR21 U316 ( .A(n35), .B(n82), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [8]) );
  INV3 U317 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[6][1] ), .Q(n82) );
  INV3 U318 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[5][5] ), .Q(n192) );
  INV3 U319 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[5][5] ), .Q(n182) );
  INV3 U320 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[5][5] ), .Q(n170) );
  INV3 U321 ( .A(n223), .Q(n193) );
  NAND22 U322 ( .A(\send_ppm1/dp_cluster_4/mult_123/A2[8] ), .B(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[5][5] ), .Q(n223) );
  INV3 U323 ( .A(n229), .Q(n183) );
  NAND22 U324 ( .A(\send_ppm1/dp_cluster_3/mult_120/A2[8] ), .B(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[5][5] ), .Q(n229) );
  INV3 U325 ( .A(n235), .Q(n171) );
  NAND22 U326 ( .A(\send_ppm1/dp_cluster_2/mult_117/A2[8] ), .B(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[5][5] ), .Q(n235) );
  NOR21 U327 ( .A(n147), .B(n244), .Q(n243) );
  NAND22 U328 ( .A(n151), .B(\send_ppm1/dp_cluster_1/mult_114/SUMB[6][5] ), 
        .Q(n244) );
  NOR21 U329 ( .A(n189), .B(n226), .Q(n225) );
  NAND22 U330 ( .A(n193), .B(\send_ppm1/dp_cluster_4/mult_123/SUMB[6][5] ), 
        .Q(n226) );
  NOR21 U331 ( .A(n181), .B(n232), .Q(n231) );
  NAND22 U332 ( .A(n183), .B(\send_ppm1/dp_cluster_3/mult_120/SUMB[6][5] ), 
        .Q(n232) );
  NOR21 U333 ( .A(n167), .B(n238), .Q(n237) );
  NAND22 U334 ( .A(n171), .B(\send_ppm1/dp_cluster_2/mult_117/SUMB[6][5] ), 
        .Q(n238) );
  INV3 U335 ( .A(n32), .Q(\send_ppm1/sig_cyclesTrame1 [15]) );
  NOR21 U336 ( .A(\send_ppm1/dp_cluster_1/N263 ), .B(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [14]), .Q(n32) );
  INV3 U337 ( .A(n45), .Q(\send_ppm1/dp_cluster_4/sub_123_cf/carry [7]) );
  NOR21 U338 ( .A(\send_ppm1/dp_cluster_4/mult_123/SUMB[5][1] ), .B(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [6]), .Q(n45) );
  INV3 U339 ( .A(n40), .Q(\send_ppm1/dp_cluster_3/sub_120_cf/carry [7]) );
  NOR21 U340 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[5][1] ), .B(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [6]), .Q(n40) );
  INV3 U341 ( .A(n35), .Q(\send_ppm1/dp_cluster_2/sub_117_cf/carry [7]) );
  NOR21 U342 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[5][1] ), .B(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [6]), .Q(n35) );
  INV3 U343 ( .A(\send_ppm1/dp_cluster_1/mult_114/CARRYB[7][5] ), .Q(n66) );
  NOR21 U344 ( .A(n92), .B(n93), .Q(\send_ppm1/dp_cluster_3/mult_120/A2[8] )
         );
  INV3 U345 ( .A(\send_ppm1/dp_cluster_3/mult_120/CARRYB[7][1] ), .Q(n92) );
  INV3 U346 ( .A(\send_ppm1/dp_cluster_3/mult_120/SUMB[4][5] ), .Q(n93) );
  NOR21 U347 ( .A(n78), .B(n79), .Q(\send_ppm1/dp_cluster_2/mult_117/A2[8] )
         );
  INV3 U348 ( .A(\send_ppm1/dp_cluster_2/mult_117/CARRYB[7][1] ), .Q(n78) );
  INV3 U349 ( .A(\send_ppm1/dp_cluster_2/mult_117/SUMB[4][5] ), .Q(n79) );
  INV3 U350 ( .A(n37), .Q(\send_ppm1/sig_cyclesTrame2 [15]) );
  NOR21 U351 ( .A(\send_ppm1/dp_cluster_2/N248 ), .B(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [14]), .Q(n37) );
  INV3 U352 ( .A(n42), .Q(\send_ppm1/sig_cyclesTrame3 [15]) );
  NOR21 U353 ( .A(\send_ppm1/dp_cluster_3/N233 ), .B(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [14]), .Q(n42) );
  INV3 U354 ( .A(n47), .Q(\send_ppm1/sig_cyclesTrame4 [15]) );
  NOR21 U355 ( .A(\send_ppm1/dp_cluster_4/N218 ), .B(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [14]), .Q(n47) );
  INV3 U356 ( .A(\send_ppm1/dp_cluster_4/mult_123/CARRYB[7][5] ), .Q(n108) );
  INV3 U357 ( .A(\send_ppm1/dp_cluster_3/mult_120/CARRYB[7][5] ), .Q(n94) );
  INV3 U358 ( .A(\send_ppm1/dp_cluster_2/mult_117/CARRYB[7][5] ), .Q(n80) );
  NOR40 U359 ( .A(n363), .B(n362), .C(n361), .D(n360), .Q(\send_ppm1/N148 ) );
  NAND41 U360 ( .A(n160), .B(n347), .C(n346), .D(n345), .Q(n363) );
  NAND41 U361 ( .A(n351), .B(n350), .C(n349), .D(n348), .Q(n362) );
  NAND41 U362 ( .A(n355), .B(n354), .C(n353), .D(n352), .Q(n361) );
  XNR21 U363 ( .A(\send_ppm1/dp_cluster_0/N296 ), .B(n23), .Q(\send_ppm1/N179 ) );
  AOI221 U364 ( .A(n3), .B(n1), .C(n1), .D(\send_ppm1/N179 ), .Q(n262) );
  NOR21 U365 ( .A(n3), .B(n13), .Q(n298) );
  NOR21 U366 ( .A(n3), .B(n14), .Q(n320) );
  INV3 U367 ( .A(n342), .Q(n160) );
  NOR21 U368 ( .A(n3), .B(n9), .Q(n342) );
  NOR21 U369 ( .A(n3), .B(n22), .Q(n276) );
  NOR31 U370 ( .A(\send_ppm1/n71 ), .B(\send_ppm1/n72 ), .C(\send_ppm1/n70 ), 
        .Q(\send_ppm1/n69 ) );
  INV3 U371 ( .A(\send_ppm1/n71 ), .Q(n203) );
  INV3 U372 ( .A(\send_ppm1/n72 ), .Q(n137) );
  INV3 U373 ( .A(\send_ppm1/n76 ), .Q(n140) );
  INV3 U374 ( .A(\send_ppm1/n60 ), .Q(n138) );
  INV3 U375 ( .A(\send_ppm1/n70 ), .Q(n132) );
  BUF2 U376 ( .A(sig_reg[28]), .Q(n123) );
  NOR21 U377 ( .A(n135), .B(n134), .Q(sig_reg[28]) );
  NAND22 U378 ( .A(n135), .B(n134), .Q(sig_reg[7]) );
  XOR21 U379 ( .A(\send_ppm1/sig_reg_storage [0]), .B(
        \send_ppm1/sig_reg_storage [1]), .Q(\send_ppm1/sig_cyclesTrame1 [2])
         );
  INV3 U380 ( .A(\send_ppm1/n73 ), .Q(n130) );
  OAI2111 U381 ( .A(n203), .B(\send_ppm1/n70 ), .C(\send_ppm1/n74 ), .D(
        \send_ppm1/n75 ), .Q(\send_ppm1/n73 ) );
  NAND31 U382 ( .A(\send_ppm1/n63 ), .B(\send_ppm1/n53 ), .C(i_reset_n_top), 
        .Q(\send_ppm1/n75 ) );
  NAND31 U383 ( .A(\send_ppm1/n76 ), .B(n141), .C(i_reset_n_top), .Q(
        \send_ppm1/n74 ) );
  XNR21 U384 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [3]), .B(
        \send_ppm1/sig_reg_storage [2]), .Q(\send_ppm1/sig_cyclesTrame1 [3])
         );
  XNR21 U385 ( .A(\send_ppm1/dp_cluster_1/sub_114_cf/carry [4]), .B(
        \send_ppm1/sig_reg_storage [3]), .Q(\send_ppm1/sig_cyclesTrame1 [4])
         );
  NAND22 U386 ( .A(\send_ppm1/sig_state [0]), .B(\send_ppm1/n58 ), .Q(
        \send_ppm1/n65 ) );
  INV3 U387 ( .A(\send_ppm1/n69 ), .Q(n133) );
  INV3 U388 ( .A(\send_ppm1/n66 ), .Q(n129) );
  NOR21 U389 ( .A(n9), .B(n6), .Q(\send_ppm1/dp_cluster_1/sub_114_cf/carry [3]) );
  NOR21 U390 ( .A(\send_ppm1/dp_cluster_1/mult_114/SUMB[1][5] ), .B(n9), .Q(
        \send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [3]) );
  NAND41 U391 ( .A(\send_ppm1/n69 ), .B(\send_ppm1/sig_state [1]), .C(
        \send_ppm1/sig_state [0]), .D(\send_ppm1/n57 ), .Q(\send_ppm1/n68 ) );
  AOI211 U392 ( .A(n132), .B(\send_ppm1/n58 ), .C(\send_ppm1/n66 ), .Q(
        \send_ppm1/n67 ) );
  XNR21 U393 ( .A(\send_ppm1/N194 ), .B(\send_ppm1/sig_out_local_count [16]), 
        .Q(n252) );
  INV3 U394 ( .A(n48), .Q(
        \send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [2]) );
  INV3 U395 ( .A(\send_ppm1/sig_cyclesTrame4 [2]), .Q(n201) );
  XOR21 U396 ( .A(\send_ppm1/sig_reg_storage [0]), .B(n159), .Q(
        \send_ppm1/dp_cluster_0/N18 ) );
  NAND22 U397 ( .A(i_reset_n_top), .B(n136), .Q(\send_ppm1/local_counter1/n22 ) );
  INV3 U398 ( .A(\send_ppm1/sig_in_init ), .Q(n136) );
  OAI2111 U399 ( .A(n140), .B(n141), .C(\send_ppm1/n60 ), .D(\send_ppm1/n61 ), 
        .Q(\send_ppm1/sig_in_init ) );
  AOI221 U400 ( .A(n203), .B(\send_ppm1/n62 ), .C(\send_ppm1/n63 ), .D(
        \send_ppm1/n64 ), .Q(\send_ppm1/n61 ) );
  XNR21 U401 ( .A(\send_ppm1/N197 ), .B(\send_ppm1/sig_out_local_count [19]), 
        .Q(n266) );
  XNR21 U402 ( .A(\send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [19]), 
        .B(\send_ppm1/dp_cluster_0/N278 ), .Q(\send_ppm1/N197 ) );
  XNR21 U403 ( .A(\send_ppm1/dp_cluster_0/add_1_root_sub_235_cf/carry [19]), 
        .B(\send_ppm1/dp_cluster_0/sub_4_root_sub_235_cf/carry [16]), .Q(
        \send_ppm1/dp_cluster_0/N278 ) );
  INV3 U404 ( .A(n55), .Q(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [19]) );
  INV3 U405 ( .A(n28), .Q(\send_ppm1/dp_cluster_1/sub_114_cf/carry [4]) );
  NOR21 U406 ( .A(\send_ppm1/sig_reg_storage [2]), .B(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [3]), .Q(n28) );
  NAND22 U407 ( .A(n256), .B(n255), .Q(n257) );
  XNR21 U408 ( .A(\send_ppm1/N195 ), .B(\send_ppm1/sig_out_local_count [17]), 
        .Q(n255) );
  XNR21 U409 ( .A(\send_ppm1/N196 ), .B(\send_ppm1/sig_out_local_count [18]), 
        .Q(n256) );
  XNR21 U410 ( .A(\send_ppm1/dp_cluster_0/N280 ), .B(
        \send_ppm1/dp_cluster_0/sub_0_root_sub_235_cf/carry [17]), .Q(
        \send_ppm1/N195 ) );
  NOR21 U411 ( .A(n120), .B(\send_ppm1/local_counter1/v_val [0]), .Q(
        \send_ppm1/local_counter1/N46 ) );
  XNR21 U412 ( .A(\send_ppm1/local_counter1/add_34/carry [19]), .B(
        \send_ppm1/local_counter1/v_val [19]), .Q(n24) );
  XOR21 U413 ( .A(\send_ppm1/sig_reg_storage [8]), .B(
        \send_ppm1/sig_reg_storage [9]), .Q(\send_ppm1/sig_cyclesTrame2 [2])
         );
  XOR21 U414 ( .A(\send_ppm1/sig_reg_storage [16]), .B(
        \send_ppm1/sig_reg_storage [17]), .Q(\send_ppm1/sig_cyclesTrame3 [2])
         );
  XNR21 U415 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [3]), .B(
        \send_ppm1/sig_reg_storage [10]), .Q(\send_ppm1/sig_cyclesTrame2 [3])
         );
  XNR21 U416 ( .A(\send_ppm1/dp_cluster_2/sub_117_cf/carry [4]), .B(
        \send_ppm1/sig_reg_storage [11]), .Q(\send_ppm1/sig_cyclesTrame2 [4])
         );
  XNR21 U417 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [3]), .B(
        \send_ppm1/sig_reg_storage [18]), .Q(\send_ppm1/sig_cyclesTrame3 [3])
         );
  XNR21 U418 ( .A(\send_ppm1/dp_cluster_3/sub_120_cf/carry [4]), .B(
        \send_ppm1/sig_reg_storage [19]), .Q(\send_ppm1/sig_cyclesTrame3 [4])
         );
  XOR21 U419 ( .A(\send_ppm1/sig_reg_storage [24]), .B(
        \send_ppm1/sig_reg_storage [25]), .Q(\send_ppm1/sig_cyclesTrame4 [2])
         );
  XOR21 U420 ( .A(\send_ppm1/sig_reg_storage [4]), .B(
        \send_ppm1/sig_reg_storage [0]), .Q(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[4][1] ) );
  XNR21 U421 ( .A(n242), .B(\send_ppm1/dp_cluster_1/mult_114/A2[12] ), .Q(
        \send_ppm1/dp_cluster_1/N263 ) );
  NOR21 U422 ( .A(n66), .B(n18), .Q(\send_ppm1/dp_cluster_1/mult_114/A2[12] )
         );
  NAND22 U423 ( .A(\send_ppm1/dp_cluster_1/mult_114/A1[11] ), .B(n243), .Q(
        n242) );
  XNR21 U424 ( .A(n9), .B(\send_ppm1/sig_reg_storage [24]), .Q(
        \send_ppm1/dp_cluster_0/N296 ) );
  XOR21 U425 ( .A(\send_ppm1/sig_reg_storage [7]), .B(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[7][5] ), .Q(
        \send_ppm1/dp_cluster_1/mult_114/A1[11] ) );
  XNR21 U426 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [3]), .B(
        \send_ppm1/sig_reg_storage [26]), .Q(\send_ppm1/sig_cyclesTrame4 [3])
         );
  XNR21 U427 ( .A(\send_ppm1/dp_cluster_4/sub_123_cf/carry [4]), .B(
        \send_ppm1/sig_reg_storage [27]), .Q(\send_ppm1/sig_cyclesTrame4 [4])
         );
  NOR21 U428 ( .A(\send_ppm1/sig_reg_storage [24]), .B(n9), .Q(n48) );
  NOR21 U429 ( .A(n22), .B(n15), .Q(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [3]) );
  NOR21 U430 ( .A(n22), .B(n15), .Q(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[1][5] ) );
  NOR21 U431 ( .A(n9), .B(n6), .Q(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[1][5] ) );
  NOR21 U432 ( .A(n7), .B(n22), .Q(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[4][1] ) );
  XOR21 U433 ( .A(\send_ppm1/sig_reg_storage [24]), .B(
        \send_ppm1/sig_reg_storage [25]), .Q(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[1][5] ) );
  NOR21 U434 ( .A(n4), .B(n9), .Q(
        \send_ppm1/dp_cluster_1/mult_114/CARRYB[4][1] ) );
  XOR21 U435 ( .A(\send_ppm1/sig_reg_storage [0]), .B(
        \send_ppm1/sig_reg_storage [1]), .Q(
        \send_ppm1/dp_cluster_1/mult_114/SUMB[1][5] ) );
  NOR21 U436 ( .A(n13), .B(n16), .Q(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[1][5] ) );
  NOR21 U437 ( .A(n14), .B(n17), .Q(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[1][5] ) );
  NOR21 U438 ( .A(n2), .B(n13), .Q(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[4][1] ) );
  XOR21 U439 ( .A(\send_ppm1/sig_reg_storage [16]), .B(
        \send_ppm1/sig_reg_storage [17]), .Q(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[1][5] ) );
  NOR21 U440 ( .A(n13), .B(n16), .Q(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [3]) );
  NOR21 U441 ( .A(n14), .B(n17), .Q(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [3]) );
  XNR21 U442 ( .A(\send_ppm1/N193 ), .B(\send_ppm1/sig_out_local_count [15]), 
        .Q(n254) );
  INV3 U443 ( .A(n43), .Q(\send_ppm1/dp_cluster_4/sub_123_cf/carry [4]) );
  NOR21 U444 ( .A(\send_ppm1/sig_reg_storage [26]), .B(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [3]), .Q(n43) );
  INV3 U445 ( .A(n38), .Q(\send_ppm1/dp_cluster_3/sub_120_cf/carry [4]) );
  NOR21 U446 ( .A(\send_ppm1/sig_reg_storage [18]), .B(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [3]), .Q(n38) );
  INV3 U447 ( .A(n33), .Q(\send_ppm1/dp_cluster_2/sub_117_cf/carry [4]) );
  NOR21 U448 ( .A(\send_ppm1/sig_reg_storage [10]), .B(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [3]), .Q(n33) );
  INV3 U449 ( .A(n29), .Q(\send_ppm1/dp_cluster_1/sub_114_cf/carry [5]) );
  NOR21 U450 ( .A(\send_ppm1/sig_reg_storage [3]), .B(
        \send_ppm1/dp_cluster_1/sub_114_cf/carry [4]), .Q(n29) );
  INV3 U451 ( .A(n44), .Q(\send_ppm1/dp_cluster_4/sub_123_cf/carry [5]) );
  NOR21 U452 ( .A(\send_ppm1/sig_reg_storage [27]), .B(
        \send_ppm1/dp_cluster_4/sub_123_cf/carry [4]), .Q(n44) );
  INV3 U453 ( .A(n39), .Q(\send_ppm1/dp_cluster_3/sub_120_cf/carry [5]) );
  NOR21 U454 ( .A(\send_ppm1/sig_reg_storage [19]), .B(
        \send_ppm1/dp_cluster_3/sub_120_cf/carry [4]), .Q(n39) );
  INV3 U455 ( .A(n34), .Q(\send_ppm1/dp_cluster_2/sub_117_cf/carry [5]) );
  NOR21 U456 ( .A(\send_ppm1/sig_reg_storage [11]), .B(
        \send_ppm1/dp_cluster_2/sub_117_cf/carry [4]), .Q(n34) );
  INV3 U457 ( .A(\send_ppm1/n77 ), .Q(n131) );
  NAND31 U458 ( .A(i_reset_n_top), .B(\send_ppm1/n76 ), .C(\send_ppm1/N198 ), 
        .Q(\send_ppm1/n77 ) );
  XOR21 U459 ( .A(\send_ppm1/sig_reg_storage [28]), .B(
        \send_ppm1/sig_reg_storage [24]), .Q(
        \send_ppm1/dp_cluster_4/mult_123/SUMB[4][1] ) );
  XOR21 U460 ( .A(\send_ppm1/sig_reg_storage [20]), .B(
        \send_ppm1/sig_reg_storage [16]), .Q(
        \send_ppm1/dp_cluster_3/mult_120/SUMB[4][1] ) );
  XOR21 U461 ( .A(\send_ppm1/sig_reg_storage [12]), .B(
        \send_ppm1/sig_reg_storage [8]), .Q(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[4][1] ) );
  XNR21 U462 ( .A(n224), .B(\send_ppm1/dp_cluster_4/mult_123/A2[12] ), .Q(
        \send_ppm1/dp_cluster_4/N218 ) );
  NOR21 U463 ( .A(n108), .B(n19), .Q(\send_ppm1/dp_cluster_4/mult_123/A2[12] )
         );
  NAND22 U464 ( .A(\send_ppm1/dp_cluster_4/mult_123/A1[11] ), .B(n225), .Q(
        n224) );
  XNR21 U465 ( .A(n236), .B(\send_ppm1/dp_cluster_2/mult_117/A2[12] ), .Q(
        \send_ppm1/dp_cluster_2/N248 ) );
  NOR21 U466 ( .A(n80), .B(n20), .Q(\send_ppm1/dp_cluster_2/mult_117/A2[12] )
         );
  NAND22 U467 ( .A(\send_ppm1/dp_cluster_2/mult_117/A1[11] ), .B(n237), .Q(
        n236) );
  XOR21 U468 ( .A(\send_ppm1/sig_reg_storage [31]), .B(
        \send_ppm1/dp_cluster_4/mult_123/CARRYB[7][5] ), .Q(
        \send_ppm1/dp_cluster_4/mult_123/A1[11] ) );
  XOR21 U469 ( .A(\send_ppm1/sig_reg_storage [23]), .B(
        \send_ppm1/dp_cluster_3/mult_120/CARRYB[7][5] ), .Q(
        \send_ppm1/dp_cluster_3/mult_120/A1[11] ) );
  XOR21 U470 ( .A(\send_ppm1/sig_reg_storage [15]), .B(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[7][5] ), .Q(
        \send_ppm1/dp_cluster_2/mult_117/A1[11] ) );
  OAI2111 U471 ( .A(\send_ppm1/N198 ), .B(n140), .C(\send_ppm1/n78 ), .D(
        i_reset_n_top), .Q(\send_ppm1/N82 ) );
  NAND31 U472 ( .A(\send_ppm1/n72 ), .B(n203), .C(\send_ppm1/n79 ), .Q(
        \send_ppm1/n78 ) );
  NOR21 U473 ( .A(n8), .B(n14), .Q(
        \send_ppm1/dp_cluster_2/mult_117/CARRYB[4][1] ) );
  XOR21 U474 ( .A(\send_ppm1/sig_reg_storage [8]), .B(
        \send_ppm1/sig_reg_storage [9]), .Q(
        \send_ppm1/dp_cluster_2/mult_117/SUMB[1][5] ) );
  XNR21 U475 ( .A(\send_ppm1/N192 ), .B(\send_ppm1/sig_out_local_count [14]), 
        .Q(n253) );
  XNR21 U476 ( .A(n230), .B(\send_ppm1/dp_cluster_3/mult_120/A2[12] ), .Q(
        \send_ppm1/dp_cluster_3/N233 ) );
  NOR21 U477 ( .A(n94), .B(n21), .Q(\send_ppm1/dp_cluster_3/mult_120/A2[12] )
         );
  NAND22 U478 ( .A(\send_ppm1/dp_cluster_3/mult_120/A1[11] ), .B(n231), .Q(
        n230) );
  XNR21 U479 ( .A(\send_ppm1/N190 ), .B(\send_ppm1/sig_out_local_count [12]), 
        .Q(n250) );
  XNR21 U480 ( .A(\send_ppm1/N191 ), .B(\send_ppm1/sig_out_local_count [13]), 
        .Q(n251) );
  XNR21 U481 ( .A(\send_ppm1/N189 ), .B(\send_ppm1/sig_out_local_count [11]), 
        .Q(n247) );
  XNR21 U482 ( .A(\send_ppm1/N188 ), .B(\send_ppm1/sig_out_local_count [10]), 
        .Q(n249) );
  XNR21 U483 ( .A(\send_ppm1/N187 ), .B(\send_ppm1/sig_out_local_count [9]), 
        .Q(n248) );
  NAND41 U484 ( .A(n334), .B(n337), .C(n336), .D(n335), .Q(n338) );
  NOR40 U485 ( .A(\send_ppm1/sig_out_local_count [19]), .B(
        \send_ppm1/sig_out_local_count [18]), .C(
        \send_ppm1/sig_out_local_count [17]), .D(
        \send_ppm1/sig_out_local_count [16]), .Q(n334) );
  XNR21 U486 ( .A(\send_ppm1/sig_cyclesTrame2 [13]), .B(
        \send_ppm1/sig_out_local_count [13]), .Q(n335) );
  XNR21 U487 ( .A(\send_ppm1/sig_cyclesTrame2 [15]), .B(
        \send_ppm1/sig_out_local_count [15]), .Q(n337) );
  NAND41 U488 ( .A(n312), .B(n315), .C(n314), .D(n313), .Q(n316) );
  NOR40 U489 ( .A(\send_ppm1/sig_out_local_count [19]), .B(
        \send_ppm1/sig_out_local_count [18]), .C(
        \send_ppm1/sig_out_local_count [17]), .D(
        \send_ppm1/sig_out_local_count [16]), .Q(n312) );
  XNR21 U490 ( .A(\send_ppm1/sig_cyclesTrame3 [13]), .B(
        \send_ppm1/sig_out_local_count [13]), .Q(n313) );
  XNR21 U491 ( .A(\send_ppm1/sig_cyclesTrame3 [15]), .B(
        \send_ppm1/sig_out_local_count [15]), .Q(n315) );
  NAND41 U492 ( .A(n356), .B(n359), .C(n358), .D(n357), .Q(n360) );
  NOR40 U493 ( .A(\send_ppm1/sig_out_local_count [19]), .B(
        \send_ppm1/sig_out_local_count [18]), .C(
        \send_ppm1/sig_out_local_count [17]), .D(
        \send_ppm1/sig_out_local_count [16]), .Q(n356) );
  XNR21 U494 ( .A(\send_ppm1/sig_cyclesTrame1 [13]), .B(
        \send_ppm1/sig_out_local_count [13]), .Q(n357) );
  XNR21 U495 ( .A(\send_ppm1/sig_cyclesTrame1 [15]), .B(
        \send_ppm1/sig_out_local_count [15]), .Q(n359) );
  INV3 U496 ( .A(\send_ppm1/N169 ), .Q(n185) );
  AOI311 U497 ( .A(\send_ppm1/N148 ), .B(\send_ppm1/n58 ), .C(
        \send_ppm1/sig_state [0]), .D(\send_ppm1/n92 ), .Q(\send_ppm1/n91 ) );
  NOR40 U498 ( .A(n297), .B(n296), .C(n295), .D(n294), .Q(\send_ppm1/N169 ) );
  XNR21 U499 ( .A(\send_ppm1/sig_cyclesTrame2 [14]), .B(
        \send_ppm1/sig_out_local_count [14]), .Q(n336) );
  XNR21 U500 ( .A(\send_ppm1/sig_cyclesTrame3 [14]), .B(
        \send_ppm1/sig_out_local_count [14]), .Q(n314) );
  XNR21 U501 ( .A(\send_ppm1/sig_cyclesTrame1 [14]), .B(
        \send_ppm1/sig_out_local_count [14]), .Q(n358) );
  NOR21 U502 ( .A(\send_ppm1/n93 ), .B(\send_ppm1/n58 ), .Q(\send_ppm1/n92 )
         );
  AOI221 U503 ( .A(\send_ppm1/N156 ), .B(\send_ppm1/n59 ), .C(\send_ppm1/N163 ), .D(\send_ppm1/sig_state [0]), .Q(\send_ppm1/n93 ) );
  NOR40 U504 ( .A(n319), .B(n318), .C(n317), .D(n316), .Q(\send_ppm1/N163 ) );
  NOR40 U505 ( .A(n341), .B(n340), .C(n339), .D(n338), .Q(\send_ppm1/N156 ) );
  NAND41 U506 ( .A(n290), .B(n293), .C(n292), .D(n291), .Q(n294) );
  NOR40 U507 ( .A(\send_ppm1/sig_out_local_count [19]), .B(
        \send_ppm1/sig_out_local_count [18]), .C(
        \send_ppm1/sig_out_local_count [17]), .D(
        \send_ppm1/sig_out_local_count [16]), .Q(n290) );
  XNR21 U508 ( .A(\send_ppm1/sig_cyclesTrame4 [13]), .B(
        \send_ppm1/sig_out_local_count [13]), .Q(n291) );
  XNR21 U509 ( .A(\send_ppm1/sig_cyclesTrame4 [15]), .B(
        \send_ppm1/sig_out_local_count [15]), .Q(n293) );
  NAND41 U510 ( .A(n333), .B(n332), .C(n331), .D(n330), .Q(n339) );
  XNR21 U511 ( .A(\send_ppm1/sig_cyclesTrame2 [9]), .B(
        \send_ppm1/sig_out_local_count [9]), .Q(n330) );
  XNR21 U512 ( .A(\send_ppm1/sig_cyclesTrame2 [10]), .B(
        \send_ppm1/sig_out_local_count [10]), .Q(n331) );
  XNR21 U513 ( .A(\send_ppm1/sig_cyclesTrame2 [11]), .B(
        \send_ppm1/sig_out_local_count [11]), .Q(n332) );
  NAND41 U514 ( .A(n311), .B(n310), .C(n309), .D(n308), .Q(n317) );
  XNR21 U515 ( .A(\send_ppm1/sig_cyclesTrame3 [9]), .B(
        \send_ppm1/sig_out_local_count [9]), .Q(n308) );
  XNR21 U516 ( .A(\send_ppm1/sig_cyclesTrame3 [10]), .B(
        \send_ppm1/sig_out_local_count [10]), .Q(n309) );
  XNR21 U517 ( .A(\send_ppm1/sig_cyclesTrame3 [11]), .B(
        \send_ppm1/sig_out_local_count [11]), .Q(n310) );
  NAND41 U518 ( .A(n289), .B(n288), .C(n287), .D(n286), .Q(n295) );
  XNR21 U519 ( .A(\send_ppm1/sig_cyclesTrame4 [9]), .B(
        \send_ppm1/sig_out_local_count [9]), .Q(n286) );
  XNR21 U520 ( .A(\send_ppm1/sig_cyclesTrame4 [10]), .B(
        \send_ppm1/sig_out_local_count [10]), .Q(n287) );
  XNR21 U521 ( .A(\send_ppm1/sig_cyclesTrame4 [11]), .B(
        \send_ppm1/sig_out_local_count [11]), .Q(n288) );
  OAI2111 U522 ( .A(\send_ppm1/n64 ), .B(\send_ppm1/n80 ), .C(\send_ppm1/n81 ), 
        .D(i_reset_n_top), .Q(\send_ppm1/N81 ) );
  NAND22 U523 ( .A(\send_ppm1/n63 ), .B(\send_ppm1/n53 ), .Q(\send_ppm1/n80 )
         );
  NAND31 U524 ( .A(n203), .B(n137), .C(\send_ppm1/n79 ), .Q(\send_ppm1/n81 )
         );
  XNR21 U525 ( .A(\send_ppm1/N185 ), .B(\send_ppm1/sig_out_local_count [7]), 
        .Q(n271) );
  XNR21 U526 ( .A(\send_ppm1/sig_cyclesTrame2 [12]), .B(
        \send_ppm1/sig_out_local_count [12]), .Q(n333) );
  XNR21 U527 ( .A(\send_ppm1/sig_cyclesTrame3 [12]), .B(
        \send_ppm1/sig_out_local_count [12]), .Q(n311) );
  XNR21 U528 ( .A(\send_ppm1/sig_cyclesTrame1 [12]), .B(
        \send_ppm1/sig_out_local_count [12]), .Q(n355) );
  XNR21 U529 ( .A(\send_ppm1/sig_cyclesTrame4 [12]), .B(
        \send_ppm1/sig_out_local_count [12]), .Q(n289) );
  XNR21 U530 ( .A(\send_ppm1/N186 ), .B(\send_ppm1/sig_out_local_count [8]), 
        .Q(n272) );
  XNR21 U531 ( .A(\send_ppm1/sig_cyclesTrame4 [14]), .B(
        \send_ppm1/sig_out_local_count [14]), .Q(n292) );
  XNR21 U532 ( .A(\send_ppm1/N184 ), .B(\send_ppm1/sig_out_local_count [6]), 
        .Q(n268) );
  XNR21 U533 ( .A(\send_ppm1/sig_cyclesTrame1 [11]), .B(
        \send_ppm1/sig_out_local_count [11]), .Q(n354) );
  NAND41 U534 ( .A(n329), .B(n328), .C(n327), .D(n326), .Q(n340) );
  XNR21 U535 ( .A(\send_ppm1/sig_cyclesTrame2 [5]), .B(
        \send_ppm1/sig_out_local_count [5]), .Q(n326) );
  XNR21 U536 ( .A(\send_ppm1/sig_cyclesTrame2 [6]), .B(
        \send_ppm1/sig_out_local_count [6]), .Q(n327) );
  XNR21 U537 ( .A(\send_ppm1/sig_cyclesTrame2 [7]), .B(
        \send_ppm1/sig_out_local_count [7]), .Q(n328) );
  NAND41 U538 ( .A(n307), .B(n306), .C(n305), .D(n304), .Q(n318) );
  XNR21 U539 ( .A(\send_ppm1/sig_cyclesTrame3 [5]), .B(
        \send_ppm1/sig_out_local_count [5]), .Q(n304) );
  XNR21 U540 ( .A(\send_ppm1/sig_cyclesTrame3 [6]), .B(
        \send_ppm1/sig_out_local_count [6]), .Q(n305) );
  XNR21 U541 ( .A(\send_ppm1/sig_cyclesTrame3 [7]), .B(
        \send_ppm1/sig_out_local_count [7]), .Q(n306) );
  XNR21 U542 ( .A(\send_ppm1/sig_cyclesTrame2 [8]), .B(
        \send_ppm1/sig_out_local_count [8]), .Q(n329) );
  XNR21 U543 ( .A(\send_ppm1/sig_cyclesTrame3 [8]), .B(
        \send_ppm1/sig_out_local_count [8]), .Q(n307) );
  XNR21 U544 ( .A(\send_ppm1/N182 ), .B(\send_ppm1/sig_out_local_count [4]), 
        .Q(n269) );
  XNR21 U545 ( .A(\send_ppm1/N183 ), .B(\send_ppm1/sig_out_local_count [5]), 
        .Q(n270) );
  XNR21 U546 ( .A(\send_ppm1/sig_cyclesTrame1 [10]), .B(
        \send_ppm1/sig_out_local_count [10]), .Q(n353) );
  XNR21 U547 ( .A(\send_ppm1/sig_cyclesTrame1 [9]), .B(
        \send_ppm1/sig_out_local_count [9]), .Q(n352) );
  NAND41 U548 ( .A(n285), .B(n284), .C(n283), .D(n282), .Q(n296) );
  XNR21 U549 ( .A(\send_ppm1/sig_cyclesTrame4 [5]), .B(
        \send_ppm1/sig_out_local_count [5]), .Q(n282) );
  XNR21 U550 ( .A(\send_ppm1/sig_cyclesTrame4 [6]), .B(
        \send_ppm1/sig_out_local_count [6]), .Q(n283) );
  XNR21 U551 ( .A(\send_ppm1/sig_cyclesTrame4 [7]), .B(
        \send_ppm1/sig_out_local_count [7]), .Q(n284) );
  XOR21 U552 ( .A(\send_ppm1/N180 ), .B(\send_ppm1/sig_out_local_count [2]), 
        .Q(n264) );
  XOR21 U553 ( .A(\send_ppm1/N181 ), .B(\send_ppm1/sig_out_local_count [3]), 
        .Q(n263) );
  XNR21 U554 ( .A(\send_ppm1/sig_cyclesTrame1 [8]), .B(
        \send_ppm1/sig_out_local_count [8]), .Q(n351) );
  XNR21 U555 ( .A(\send_ppm1/sig_cyclesTrame4 [8]), .B(
        \send_ppm1/sig_out_local_count [8]), .Q(n285) );
  XNR21 U556 ( .A(\send_ppm1/sig_cyclesTrame1 [7]), .B(
        \send_ppm1/sig_out_local_count [7]), .Q(n350) );
  XNR21 U557 ( .A(\send_ppm1/sig_cyclesTrame1 [6]), .B(
        \send_ppm1/sig_out_local_count [6]), .Q(n349) );
  NAND41 U558 ( .A(n180), .B(n325), .C(n324), .D(n323), .Q(n341) );
  INV3 U559 ( .A(n320), .Q(n180) );
  XNR21 U560 ( .A(\send_ppm1/sig_cyclesTrame2 [2]), .B(
        \send_ppm1/sig_out_local_count [2]), .Q(n324) );
  NAND41 U561 ( .A(n184), .B(n303), .C(n302), .D(n301), .Q(n319) );
  INV3 U562 ( .A(n298), .Q(n184) );
  XNR21 U563 ( .A(\send_ppm1/sig_cyclesTrame3 [2]), .B(
        \send_ppm1/sig_out_local_count [2]), .Q(n302) );
  XNR21 U564 ( .A(\send_ppm1/sig_cyclesTrame1 [5]), .B(
        \send_ppm1/sig_out_local_count [5]), .Q(n348) );
  NOR21 U565 ( .A(n322), .B(n321), .Q(n323) );
  XOR21 U566 ( .A(\send_ppm1/sig_cyclesTrame2 [3]), .B(
        \send_ppm1/sig_out_local_count [3]), .Q(n322) );
  XOR21 U567 ( .A(\send_ppm1/sig_cyclesTrame2 [4]), .B(
        \send_ppm1/sig_out_local_count [4]), .Q(n321) );
  NOR21 U568 ( .A(n300), .B(n299), .Q(n301) );
  XOR21 U569 ( .A(\send_ppm1/sig_cyclesTrame3 [3]), .B(
        \send_ppm1/sig_out_local_count [3]), .Q(n300) );
  XOR21 U570 ( .A(\send_ppm1/sig_cyclesTrame3 [4]), .B(
        \send_ppm1/sig_out_local_count [4]), .Q(n299) );
  NOR21 U571 ( .A(n344), .B(n343), .Q(n345) );
  XOR21 U572 ( .A(\send_ppm1/sig_cyclesTrame1 [3]), .B(
        \send_ppm1/sig_out_local_count [3]), .Q(n344) );
  XOR21 U573 ( .A(\send_ppm1/sig_cyclesTrame1 [4]), .B(
        \send_ppm1/sig_out_local_count [4]), .Q(n343) );
  NAND41 U574 ( .A(n202), .B(n281), .C(n280), .D(n279), .Q(n297) );
  INV3 U575 ( .A(n276), .Q(n202) );
  XNR21 U576 ( .A(\send_ppm1/sig_cyclesTrame4 [2]), .B(
        \send_ppm1/sig_out_local_count [2]), .Q(n280) );
  XNR21 U577 ( .A(\send_ppm1/sig_cyclesTrame1 [2]), .B(
        \send_ppm1/sig_out_local_count [2]), .Q(n346) );
  NOR21 U578 ( .A(n278), .B(n277), .Q(n279) );
  XOR21 U579 ( .A(\send_ppm1/sig_cyclesTrame4 [3]), .B(
        \send_ppm1/sig_out_local_count [3]), .Q(n278) );
  XOR21 U580 ( .A(\send_ppm1/sig_cyclesTrame4 [4]), .B(
        \send_ppm1/sig_out_local_count [4]), .Q(n277) );
  NAND41 U581 ( .A(\send_ppm1/n82 ), .B(\send_ppm1/n83 ), .C(\send_ppm1/n84 ), 
        .D(\send_ppm1/n85 ), .Q(\send_ppm1/n71 ) );
  NOR21 U582 ( .A(\send_ppm1/sig_out_local_count [16]), .B(
        \send_ppm1/sig_out_local_count [15]), .Q(\send_ppm1/n82 ) );
  NOR31 U583 ( .A(\send_ppm1/sig_out_local_count [17]), .B(
        \send_ppm1/sig_out_local_count [19]), .C(
        \send_ppm1/sig_out_local_count [18]), .Q(\send_ppm1/n83 ) );
  NOR40 U584 ( .A(\send_ppm1/sig_out_local_count [5]), .B(n204), .C(
        \send_ppm1/sig_out_local_count [4]), .D(
        \send_ppm1/sig_out_local_count [2]), .Q(\send_ppm1/n84 ) );
  NOR31 U585 ( .A(\send_ppm1/sig_state [0]), .B(\send_ppm1/sig_state [1]), .C(
        \send_ppm1/n57 ), .Q(\send_ppm1/n72 ) );
  NOR31 U586 ( .A(\send_ppm1/n86 ), .B(\send_ppm1/n87 ), .C(\send_ppm1/n88 ), 
        .Q(\send_ppm1/n85 ) );
  NAND22 U587 ( .A(\send_ppm1/sig_out_local_count [8]), .B(
        \send_ppm1/sig_out_local_count [6]), .Q(\send_ppm1/n88 ) );
  NAND31 U588 ( .A(\send_ppm1/sig_out_local_count [1]), .B(
        \send_ppm1/sig_out_local_count [12]), .C(
        \send_ppm1/sig_out_local_count [3]), .Q(\send_ppm1/n87 ) );
  NAND41 U589 ( .A(\send_ppm1/sig_out_local_count [11]), .B(
        \send_ppm1/sig_out_local_count [10]), .C(\send_ppm1/n89 ), .D(
        \send_ppm1/sig_out_local_count [0]), .Q(\send_ppm1/n86 ) );
  NOR21 U590 ( .A(\send_ppm1/sig_out_local_count [14]), .B(
        \send_ppm1/sig_out_local_count [13]), .Q(\send_ppm1/n89 ) );
  INV3 U591 ( .A(\send_ppm1/n90 ), .Q(n204) );
  NOR21 U592 ( .A(\send_ppm1/sig_out_local_count [9]), .B(
        \send_ppm1/sig_out_local_count [7]), .Q(\send_ppm1/n90 ) );
  NOR31 U593 ( .A(\send_ppm1/current_state [0]), .B(
        \send_ppm1/current_state [2]), .C(\send_ppm1/n53 ), .Q(\send_ppm1/n76 ) );
  AOI221 U594 ( .A(\send_ppm1/n63 ), .B(\send_ppm1/current_state [1]), .C(
        \send_ppm1/n62 ), .D(\send_ppm1/current_state [2]), .Q(\send_ppm1/n60 ) );
  NAND22 U595 ( .A(i_reset_n_top), .B(\send_ppm1/n79 ), .Q(\send_ppm1/n70 ) );
  NOR21 U596 ( .A(\send_ppm1/n55 ), .B(\send_ppm1/current_state [2]), .Q(
        \send_ppm1/n63 ) );
  NOR21 U597 ( .A(\send_ppm1/current_state [0]), .B(
        \send_ppm1/current_state [1]), .Q(\send_ppm1/n62 ) );
  NOR21 U598 ( .A(n139), .B(\send_ppm1/current_state [2]), .Q(\send_ppm1/n79 )
         );
  INV3 U599 ( .A(\send_ppm1/n62 ), .Q(n139) );
  INV3 U600 ( .A(sig_reg[31]), .Q(n134) );
  INV3 U601 ( .A(sig_reg[30]), .Q(n135) );
  OAI222 U602 ( .A(n1), .B(n3), .C(n22), .D(n1), .Q(n281) );
  OAI222 U603 ( .A(n1), .B(n3), .C(n13), .D(n1), .Q(n303) );
  OAI222 U604 ( .A(n1), .B(n3), .C(n14), .D(n1), .Q(n325) );
  OAI222 U605 ( .A(n1), .B(n3), .C(n9), .D(n1), .Q(n347) );
endmodule

