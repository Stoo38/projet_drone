
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_ppm is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_top_ppm;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_ppm.all;

entity top_ppm is

   port( i_clk_top, i_reset_n_top : in std_logic;  i_sel_top : in 
         std_logic_vector (1 downto 0);  o_ppm_top : out std_logic);

end top_ppm;

architecture SYN_rtl of top_ppm is

   component OAI222
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component INV3
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND22
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI221
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND41
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR40
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI311
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI211
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component BUF2
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX22
      port( A, B, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFE1
      port( D, E, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DF3
      port( D, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component JK3
      port( J, K, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component ADD32
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADD22
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI212
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   signal sig_reg_28_port, sig_reg_7_port, send_ppm1_n95, send_ppm1_n94, 
      send_ppm1_n93, send_ppm1_n92, send_ppm1_n91, send_ppm1_n90, send_ppm1_n89
      , send_ppm1_n88, send_ppm1_n87, send_ppm1_n86, send_ppm1_n85, 
      send_ppm1_n84, send_ppm1_n83, send_ppm1_n82, send_ppm1_n81, send_ppm1_n80
      , send_ppm1_n79, send_ppm1_n78, send_ppm1_n77, send_ppm1_n76, 
      send_ppm1_n75, send_ppm1_n74, send_ppm1_n73, send_ppm1_n72, send_ppm1_n71
      , send_ppm1_n70, send_ppm1_n69, send_ppm1_n68, send_ppm1_n67, 
      send_ppm1_n66, send_ppm1_n65, send_ppm1_n64, send_ppm1_n63, send_ppm1_n62
      , send_ppm1_n61, send_ppm1_n60, send_ppm1_n59, send_ppm1_n58, 
      send_ppm1_n57, send_ppm1_n55, send_ppm1_n53, send_ppm1_dp_cluster_4_N218,
      send_ppm1_dp_cluster_4_N219, send_ppm1_dp_cluster_4_N220, 
      send_ppm1_dp_cluster_4_N221, send_ppm1_dp_cluster_4_N223, 
      send_ppm1_dp_cluster_3_N233, send_ppm1_dp_cluster_3_N234, 
      send_ppm1_dp_cluster_3_N235, send_ppm1_dp_cluster_3_N236, 
      send_ppm1_dp_cluster_3_N238, send_ppm1_dp_cluster_2_N248, 
      send_ppm1_dp_cluster_2_N249, send_ppm1_dp_cluster_2_N250, 
      send_ppm1_dp_cluster_2_N251, send_ppm1_dp_cluster_2_N253, 
      send_ppm1_dp_cluster_1_N263, send_ppm1_dp_cluster_1_N264, 
      send_ppm1_dp_cluster_1_N265, send_ppm1_dp_cluster_1_N266, 
      send_ppm1_dp_cluster_1_N268, send_ppm1_dp_cluster_0_N18, 
      send_ppm1_dp_cluster_0_N19, send_ppm1_dp_cluster_0_N20, 
      send_ppm1_dp_cluster_0_N21, send_ppm1_dp_cluster_0_N22, 
      send_ppm1_dp_cluster_0_N23, send_ppm1_dp_cluster_0_N24, 
      send_ppm1_dp_cluster_0_N25, send_ppm1_dp_cluster_0_N26, 
      send_ppm1_dp_cluster_0_N27, send_ppm1_dp_cluster_0_N278, 
      send_ppm1_dp_cluster_0_N279, send_ppm1_dp_cluster_0_N28, 
      send_ppm1_dp_cluster_0_N280, send_ppm1_dp_cluster_0_N281, 
      send_ppm1_dp_cluster_0_N282, send_ppm1_dp_cluster_0_N283, 
      send_ppm1_dp_cluster_0_N284, send_ppm1_dp_cluster_0_N285, 
      send_ppm1_dp_cluster_0_N286, send_ppm1_dp_cluster_0_N287, 
      send_ppm1_dp_cluster_0_N288, send_ppm1_dp_cluster_0_N289, 
      send_ppm1_dp_cluster_0_N29, send_ppm1_dp_cluster_0_N290, 
      send_ppm1_dp_cluster_0_N291, send_ppm1_dp_cluster_0_N292, 
      send_ppm1_dp_cluster_0_N293, send_ppm1_dp_cluster_0_N294, 
      send_ppm1_dp_cluster_0_N295, send_ppm1_dp_cluster_0_N296, 
      send_ppm1_dp_cluster_0_N30, send_ppm1_dp_cluster_0_N31, 
      send_ppm1_dp_cluster_0_N38, send_ppm1_dp_cluster_0_N39, 
      send_ppm1_dp_cluster_0_N40, send_ppm1_dp_cluster_0_N41, 
      send_ppm1_dp_cluster_0_N42, send_ppm1_dp_cluster_0_N43, 
      send_ppm1_dp_cluster_0_N44, send_ppm1_dp_cluster_0_N45, 
      send_ppm1_dp_cluster_0_N46, send_ppm1_dp_cluster_0_N47, 
      send_ppm1_dp_cluster_0_N48, send_ppm1_dp_cluster_0_N49, 
      send_ppm1_dp_cluster_0_N50, send_ppm1_dp_cluster_0_N51, send_ppm1_N198, 
      send_ppm1_N197, send_ppm1_N196, send_ppm1_N195, send_ppm1_N194, 
      send_ppm1_N193, send_ppm1_N192, send_ppm1_N191, send_ppm1_N190, 
      send_ppm1_N189, send_ppm1_N188, send_ppm1_N187, send_ppm1_N186, 
      send_ppm1_N185, send_ppm1_N184, send_ppm1_N183, send_ppm1_N182, 
      send_ppm1_N181, send_ppm1_N180, send_ppm1_N179, send_ppm1_N169, 
      send_ppm1_N163, send_ppm1_N156, send_ppm1_N148, send_ppm1_N82_port, 
      send_ppm1_N81_port, send_ppm1_sig_state_0_port, 
      send_ppm1_sig_state_1_port, send_ppm1_sig_state_2_port, 
      send_ppm1_current_state_0_port, send_ppm1_current_state_1_port, 
      send_ppm1_current_state_2_port, send_ppm1_sig_cyclesTrame4_2_port, 
      send_ppm1_sig_cyclesTrame4_3_port, send_ppm1_sig_cyclesTrame4_4_port, 
      send_ppm1_sig_cyclesTrame4_5_port, send_ppm1_sig_cyclesTrame4_6_port, 
      send_ppm1_sig_cyclesTrame4_7_port, send_ppm1_sig_cyclesTrame4_8_port, 
      send_ppm1_sig_cyclesTrame4_9_port, send_ppm1_sig_cyclesTrame4_10_port, 
      send_ppm1_sig_cyclesTrame4_11_port, send_ppm1_sig_cyclesTrame4_12_port, 
      send_ppm1_sig_cyclesTrame4_13_port, send_ppm1_sig_cyclesTrame4_14_port, 
      send_ppm1_sig_cyclesTrame4_15_port, send_ppm1_sig_cyclesTrame3_2_port, 
      send_ppm1_sig_cyclesTrame3_3_port, send_ppm1_sig_cyclesTrame3_4_port, 
      send_ppm1_sig_cyclesTrame3_5_port, send_ppm1_sig_cyclesTrame3_6_port, 
      send_ppm1_sig_cyclesTrame3_7_port, send_ppm1_sig_cyclesTrame3_8_port, 
      send_ppm1_sig_cyclesTrame3_9_port, send_ppm1_sig_cyclesTrame3_10_port, 
      send_ppm1_sig_cyclesTrame3_11_port, send_ppm1_sig_cyclesTrame3_12_port, 
      send_ppm1_sig_cyclesTrame3_13_port, send_ppm1_sig_cyclesTrame3_14_port, 
      send_ppm1_sig_cyclesTrame3_15_port, send_ppm1_sig_cyclesTrame2_2_port, 
      send_ppm1_sig_cyclesTrame2_3_port, send_ppm1_sig_cyclesTrame2_4_port, 
      send_ppm1_sig_cyclesTrame2_5_port, send_ppm1_sig_cyclesTrame2_6_port, 
      send_ppm1_sig_cyclesTrame2_7_port, send_ppm1_sig_cyclesTrame2_8_port, 
      send_ppm1_sig_cyclesTrame2_9_port, send_ppm1_sig_cyclesTrame2_10_port, 
      send_ppm1_sig_cyclesTrame2_11_port, send_ppm1_sig_cyclesTrame2_12_port, 
      send_ppm1_sig_cyclesTrame2_13_port, send_ppm1_sig_cyclesTrame2_14_port, 
      send_ppm1_sig_cyclesTrame2_15_port, send_ppm1_sig_cyclesTrame1_2_port, 
      send_ppm1_sig_cyclesTrame1_3_port, send_ppm1_sig_cyclesTrame1_4_port, 
      send_ppm1_sig_cyclesTrame1_5_port, send_ppm1_sig_cyclesTrame1_6_port, 
      send_ppm1_sig_cyclesTrame1_7_port, send_ppm1_sig_cyclesTrame1_8_port, 
      send_ppm1_sig_cyclesTrame1_9_port, send_ppm1_sig_cyclesTrame1_10_port, 
      send_ppm1_sig_cyclesTrame1_11_port, send_ppm1_sig_cyclesTrame1_12_port, 
      send_ppm1_sig_cyclesTrame1_13_port, send_ppm1_sig_cyclesTrame1_14_port, 
      send_ppm1_sig_cyclesTrame1_15_port, send_ppm1_sig_reg_storage_0_port, 
      send_ppm1_sig_reg_storage_1_port, send_ppm1_sig_reg_storage_2_port, 
      send_ppm1_sig_reg_storage_3_port, send_ppm1_sig_reg_storage_4_port, 
      send_ppm1_sig_reg_storage_5_port, send_ppm1_sig_reg_storage_6_port, 
      send_ppm1_sig_reg_storage_7_port, send_ppm1_sig_reg_storage_8_port, 
      send_ppm1_sig_reg_storage_9_port, send_ppm1_sig_reg_storage_10_port, 
      send_ppm1_sig_reg_storage_11_port, send_ppm1_sig_reg_storage_12_port, 
      send_ppm1_sig_reg_storage_13_port, send_ppm1_sig_reg_storage_14_port, 
      send_ppm1_sig_reg_storage_15_port, send_ppm1_sig_reg_storage_16_port, 
      send_ppm1_sig_reg_storage_17_port, send_ppm1_sig_reg_storage_18_port, 
      send_ppm1_sig_reg_storage_19_port, send_ppm1_sig_reg_storage_20_port, 
      send_ppm1_sig_reg_storage_21_port, send_ppm1_sig_reg_storage_22_port, 
      send_ppm1_sig_reg_storage_23_port, send_ppm1_sig_reg_storage_24_port, 
      send_ppm1_sig_reg_storage_25_port, send_ppm1_sig_reg_storage_26_port, 
      send_ppm1_sig_reg_storage_27_port, send_ppm1_sig_reg_storage_28_port, 
      send_ppm1_sig_reg_storage_29_port, send_ppm1_sig_reg_storage_30_port, 
      send_ppm1_sig_reg_storage_31_port, send_ppm1_sig_out_local_count_0_port, 
      send_ppm1_sig_out_local_count_1_port, 
      send_ppm1_sig_out_local_count_2_port, 
      send_ppm1_sig_out_local_count_3_port, 
      send_ppm1_sig_out_local_count_4_port, 
      send_ppm1_sig_out_local_count_5_port, 
      send_ppm1_sig_out_local_count_6_port, 
      send_ppm1_sig_out_local_count_7_port, 
      send_ppm1_sig_out_local_count_8_port, 
      send_ppm1_sig_out_local_count_9_port, 
      send_ppm1_sig_out_local_count_10_port, 
      send_ppm1_sig_out_local_count_11_port, 
      send_ppm1_sig_out_local_count_12_port, 
      send_ppm1_sig_out_local_count_13_port, 
      send_ppm1_sig_out_local_count_14_port, 
      send_ppm1_sig_out_local_count_15_port, 
      send_ppm1_sig_out_local_count_16_port, 
      send_ppm1_sig_out_local_count_17_port, 
      send_ppm1_sig_out_local_count_18_port, 
      send_ppm1_sig_out_local_count_19_port, send_ppm1_sig_in_init, 
      send_ppm1_local_counter1_n22, send_ppm1_local_counter1_N65, 
      send_ppm1_local_counter1_N64, send_ppm1_local_counter1_N63, 
      send_ppm1_local_counter1_N62, send_ppm1_local_counter1_N61, 
      send_ppm1_local_counter1_N60, send_ppm1_local_counter1_N59, 
      send_ppm1_local_counter1_N58, send_ppm1_local_counter1_N57, 
      send_ppm1_local_counter1_N56, send_ppm1_local_counter1_N55, 
      send_ppm1_local_counter1_N54, send_ppm1_local_counter1_N53, 
      send_ppm1_local_counter1_N52, send_ppm1_local_counter1_N51, 
      send_ppm1_local_counter1_N50, send_ppm1_local_counter1_N49, 
      send_ppm1_local_counter1_N48, send_ppm1_local_counter1_N47, 
      send_ppm1_local_counter1_N46, send_ppm1_local_counter1_N24, 
      send_ppm1_local_counter1_N23, send_ppm1_local_counter1_N22_port, 
      send_ppm1_local_counter1_N21, send_ppm1_local_counter1_N20, 
      send_ppm1_local_counter1_N19, send_ppm1_local_counter1_N18, 
      send_ppm1_local_counter1_N17, send_ppm1_local_counter1_N16, 
      send_ppm1_local_counter1_N15, send_ppm1_local_counter1_N14, 
      send_ppm1_local_counter1_N13, send_ppm1_local_counter1_N12, 
      send_ppm1_local_counter1_N11, send_ppm1_local_counter1_N10, 
      send_ppm1_local_counter1_N9, send_ppm1_local_counter1_N8, 
      send_ppm1_local_counter1_N7, send_ppm1_local_counter1_v_val_0_port, 
      send_ppm1_local_counter1_v_val_1_port, 
      send_ppm1_local_counter1_v_val_2_port, 
      send_ppm1_local_counter1_v_val_3_port, 
      send_ppm1_local_counter1_v_val_4_port, 
      send_ppm1_local_counter1_v_val_5_port, 
      send_ppm1_local_counter1_v_val_6_port, 
      send_ppm1_local_counter1_v_val_7_port, 
      send_ppm1_local_counter1_v_val_8_port, 
      send_ppm1_local_counter1_v_val_9_port, 
      send_ppm1_local_counter1_v_val_10_port, 
      send_ppm1_local_counter1_v_val_11_port, 
      send_ppm1_local_counter1_v_val_12_port, 
      send_ppm1_local_counter1_v_val_13_port, 
      send_ppm1_local_counter1_v_val_14_port, 
      send_ppm1_local_counter1_v_val_15_port, 
      send_ppm1_local_counter1_v_val_16_port, 
      send_ppm1_local_counter1_v_val_17_port, 
      send_ppm1_local_counter1_v_val_18_port, 
      send_ppm1_local_counter1_v_val_19_port, 
      send_ppm1_local_counter1_add_34_carry_2_port, 
      send_ppm1_local_counter1_add_34_carry_3_port, 
      send_ppm1_local_counter1_add_34_carry_4_port, 
      send_ppm1_local_counter1_add_34_carry_5_port, 
      send_ppm1_local_counter1_add_34_carry_6_port, 
      send_ppm1_local_counter1_add_34_carry_7_port, 
      send_ppm1_local_counter1_add_34_carry_8_port, 
      send_ppm1_local_counter1_add_34_carry_9_port, 
      send_ppm1_local_counter1_add_34_carry_10_port, 
      send_ppm1_local_counter1_add_34_carry_11_port, 
      send_ppm1_local_counter1_add_34_carry_12_port, 
      send_ppm1_local_counter1_add_34_carry_13_port, 
      send_ppm1_local_counter1_add_34_carry_14_port, 
      send_ppm1_local_counter1_add_34_carry_15_port, 
      send_ppm1_local_counter1_add_34_carry_16_port, 
      send_ppm1_local_counter1_add_34_carry_17_port, 
      send_ppm1_local_counter1_add_34_carry_18_port, 
      send_ppm1_local_counter1_add_34_carry_19_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port, 
      send_ppm1_dp_cluster_1_mult_114_A2_8_port, 
      send_ppm1_dp_cluster_1_mult_114_A2_12_port, 
      send_ppm1_dp_cluster_1_mult_114_A1_11_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port, 
      send_ppm1_dp_cluster_2_mult_117_A2_8_port, 
      send_ppm1_dp_cluster_2_mult_117_A2_12_port, 
      send_ppm1_dp_cluster_2_mult_117_A1_11_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port, 
      send_ppm1_dp_cluster_3_mult_120_A2_8_port, 
      send_ppm1_dp_cluster_3_mult_120_A2_12_port, 
      send_ppm1_dp_cluster_3_mult_120_A1_11_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port, 
      send_ppm1_dp_cluster_4_mult_123_A2_8_port, 
      send_ppm1_dp_cluster_4_mult_123_A2_12_port, 
      send_ppm1_dp_cluster_4_mult_123_A1_11_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port, n1, n2, n3, n4, n5, n6, 
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055 : std_logic;

begin
   
   send_ppm1_U39 : OAI222 port map( A => n137, B => n185, C => 
                           send_ppm1_sig_state_2_port, D => send_ppm1_n91, Q =>
                           send_ppm1_n64);
   send_ppm1_U16 : OAI212 port map( A => send_ppm1_sig_state_0_port, B => 
                           send_ppm1_n70, C => n130, Q => send_ppm1_n66);
   send_ppm1_U13 : OAI212 port map( A => send_ppm1_n67, B => send_ppm1_n57, C 
                           => send_ppm1_n68, Q => send_ppm1_n95);
   send_ppm1_U6 : OAI222 port map( A => n129, B => send_ppm1_n58, C => n133, D 
                           => send_ppm1_n65, Q => send_ppm1_n94);
   send_ppm1_local_counter1_add_34_U1_1_1 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_1_port, B => 
                           send_ppm1_local_counter1_v_val_0_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_2_port, S => 
                           send_ppm1_local_counter1_N7);
   send_ppm1_local_counter1_add_34_U1_1_2 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_2_port, B => 
                           send_ppm1_local_counter1_add_34_carry_2_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_3_port, S => 
                           send_ppm1_local_counter1_N8);
   send_ppm1_local_counter1_add_34_U1_1_3 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_3_port, B => 
                           send_ppm1_local_counter1_add_34_carry_3_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_4_port, S => 
                           send_ppm1_local_counter1_N9);
   send_ppm1_local_counter1_add_34_U1_1_4 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_4_port, B => 
                           send_ppm1_local_counter1_add_34_carry_4_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_5_port, S => 
                           send_ppm1_local_counter1_N10);
   send_ppm1_local_counter1_add_34_U1_1_5 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_5_port, B => 
                           send_ppm1_local_counter1_add_34_carry_5_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_6_port, S => 
                           send_ppm1_local_counter1_N11);
   send_ppm1_local_counter1_add_34_U1_1_6 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_6_port, B => 
                           send_ppm1_local_counter1_add_34_carry_6_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_7_port, S => 
                           send_ppm1_local_counter1_N12);
   send_ppm1_local_counter1_add_34_U1_1_7 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_7_port, B => 
                           send_ppm1_local_counter1_add_34_carry_7_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_8_port, S => 
                           send_ppm1_local_counter1_N13);
   send_ppm1_local_counter1_add_34_U1_1_8 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_8_port, B => 
                           send_ppm1_local_counter1_add_34_carry_8_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_9_port, S => 
                           send_ppm1_local_counter1_N14);
   send_ppm1_local_counter1_add_34_U1_1_9 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_9_port, B => 
                           send_ppm1_local_counter1_add_34_carry_9_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_10_port, S => 
                           send_ppm1_local_counter1_N15);
   send_ppm1_local_counter1_add_34_U1_1_10 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_10_port, B => 
                           send_ppm1_local_counter1_add_34_carry_10_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_11_port, S => 
                           send_ppm1_local_counter1_N16);
   send_ppm1_local_counter1_add_34_U1_1_11 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_11_port, B => 
                           send_ppm1_local_counter1_add_34_carry_11_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_12_port, S => 
                           send_ppm1_local_counter1_N17);
   send_ppm1_local_counter1_add_34_U1_1_12 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_12_port, B => 
                           send_ppm1_local_counter1_add_34_carry_12_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_13_port, S => 
                           send_ppm1_local_counter1_N18);
   send_ppm1_local_counter1_add_34_U1_1_13 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_13_port, B => 
                           send_ppm1_local_counter1_add_34_carry_13_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_14_port, S => 
                           send_ppm1_local_counter1_N19);
   send_ppm1_local_counter1_add_34_U1_1_14 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_14_port, B => 
                           send_ppm1_local_counter1_add_34_carry_14_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_15_port, S => 
                           send_ppm1_local_counter1_N20);
   send_ppm1_local_counter1_add_34_U1_1_15 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_15_port, B => 
                           send_ppm1_local_counter1_add_34_carry_15_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_16_port, S => 
                           send_ppm1_local_counter1_N21);
   send_ppm1_local_counter1_add_34_U1_1_16 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_16_port, B => 
                           send_ppm1_local_counter1_add_34_carry_16_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_17_port, S => 
                           send_ppm1_local_counter1_N22_port);
   send_ppm1_local_counter1_add_34_U1_1_17 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_17_port, B => 
                           send_ppm1_local_counter1_add_34_carry_17_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_18_port, S => 
                           send_ppm1_local_counter1_N23);
   send_ppm1_local_counter1_add_34_U1_1_18 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_18_port, B => 
                           send_ppm1_local_counter1_add_34_carry_18_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_19_port, S => 
                           send_ppm1_local_counter1_N24);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_2 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_2_port, B => 
                           send_ppm1_sig_cyclesTrame3_2_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_dp_cluster_0_N38);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_3 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_3_port, B => 
                           send_ppm1_sig_cyclesTrame3_3_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_dp_cluster_0_N39);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_4 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_4_port, B => 
                           send_ppm1_sig_cyclesTrame3_4_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_dp_cluster_0_N40);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_5 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_5_port, B => 
                           send_ppm1_sig_cyclesTrame3_5_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_dp_cluster_0_N41);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_6 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_6_port, B => 
                           send_ppm1_sig_cyclesTrame3_6_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_dp_cluster_0_N42);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_7 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_7_port, B => 
                           send_ppm1_sig_cyclesTrame3_7_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_dp_cluster_0_N43);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_8 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_8_port, B => 
                           send_ppm1_sig_cyclesTrame3_8_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_dp_cluster_0_N44);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_9 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_9_port, B => 
                           send_ppm1_sig_cyclesTrame3_9_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_dp_cluster_0_N45);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_10 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_10_port, B => 
                           send_ppm1_sig_cyclesTrame3_10_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_dp_cluster_0_N46);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_11 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_11_port, B => 
                           send_ppm1_sig_cyclesTrame3_11_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_dp_cluster_0_N47);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_12 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_12_port, B => 
                           send_ppm1_sig_cyclesTrame3_12_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_dp_cluster_0_N48);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_13 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_13_port, B => 
                           send_ppm1_sig_cyclesTrame3_13_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_dp_cluster_0_N49);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_14 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_14_port, B => 
                           send_ppm1_sig_cyclesTrame3_14_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_dp_cluster_0_N50);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_15 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_15_port, B => 
                           send_ppm1_sig_cyclesTrame3_15_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_dp_cluster_0_N51);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_2 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N18, B => n201, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_dp_cluster_0_N295);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_3 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N19, B => n200, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_dp_cluster_0_N294);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_4 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N20, B => n199, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_dp_cluster_0_N293);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_5 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N21, B => n198, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_dp_cluster_0_N292);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_6 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N22, B => n197, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_dp_cluster_0_N291);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_7 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N23, B => n196, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_dp_cluster_0_N290);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_8 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N24, B => n195, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_dp_cluster_0_N289);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_9 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N25, B => n194, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_dp_cluster_0_N288);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_10 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N26, B => n191, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_dp_cluster_0_N287);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_11 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N27, B => n190, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_dp_cluster_0_N286);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_12 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N28, B => n188, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_dp_cluster_0_N285);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_13 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N29, B => n187, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_dp_cluster_0_N284);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_14 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N30, B => n186, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_dp_cluster_0_N283);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_15 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N31, B => n47, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_dp_cluster_0_N282);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_2 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N295, B => n179, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_N180);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_3 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N294, B => n178, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_N181);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_4 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N293, B => n177, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_N182);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_5 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N292, B => n176, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_N183);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_6 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N291, B => n175, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_N184);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_7 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N290, B => n174, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_N185);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_8 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N289, B => n173, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_N186);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_9 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N288, B => n172, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_N187);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_10 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N287, B => n169, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_N188);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_11 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N286, B => n168, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_N189);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_12 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N285, B => n166, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_N190);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_13 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N284, B => n165, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_N191);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_14 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N283, B => n164, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_N192);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_15 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N282, B => n163, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_N193);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_16 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N281, B => n162, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, S 
                           => send_ppm1_N194);
   send_ppm1_dp_cluster_1_mult_114_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_2_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_1_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_3_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_2_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_4_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_3_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_5_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_4_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port);
   send_ppm1_dp_cluster_1_mult_114_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_5_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port);
   send_ppm1_dp_cluster_1_mult_114_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_6_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_5_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port);
   send_ppm1_dp_cluster_1_mult_114_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_6_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port);
   send_ppm1_dp_cluster_1_mult_114_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_6_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port);
   send_ppm1_dp_cluster_1_mult_114_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port);
   send_ppm1_dp_cluster_2_mult_117_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_10_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_9_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_11_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_10_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_12_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_11_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_13_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_12_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port);
   send_ppm1_dp_cluster_2_mult_117_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_13_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port);
   send_ppm1_dp_cluster_2_mult_117_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_14_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_13_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port);
   send_ppm1_dp_cluster_2_mult_117_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_14_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port);
   send_ppm1_dp_cluster_2_mult_117_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_14_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port);
   send_ppm1_dp_cluster_2_mult_117_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port);
   send_ppm1_dp_cluster_3_mult_120_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_18_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_17_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_19_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_18_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_20_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_19_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_21_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_20_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port);
   send_ppm1_dp_cluster_3_mult_120_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_21_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port);
   send_ppm1_dp_cluster_3_mult_120_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_22_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_21_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port);
   send_ppm1_dp_cluster_3_mult_120_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_22_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port);
   send_ppm1_dp_cluster_3_mult_120_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_22_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port);
   send_ppm1_dp_cluster_3_mult_120_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port);
   send_ppm1_dp_cluster_4_mult_123_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_26_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_25_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_27_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_26_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_28_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_27_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_29_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_28_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port);
   send_ppm1_dp_cluster_4_mult_123_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_29_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port);
   send_ppm1_dp_cluster_4_mult_123_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_30_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_29_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port);
   send_ppm1_dp_cluster_4_mult_123_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_30_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port);
   send_ppm1_dp_cluster_4_mult_123_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_30_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port);
   send_ppm1_dp_cluster_4_mult_123_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port);
   send_ppm1_sig_state_reg_1_inst : DF3 port map( D => send_ppm1_n94, C => 
                           i_clk_top, Q => send_ppm1_sig_state_1_port, QN => 
                           send_ppm1_n58);
   send_ppm1_current_state_reg_0_inst : DF3 port map( D => send_ppm1_N81_port, 
                           C => i_clk_top, Q => send_ppm1_current_state_0_port,
                           QN => send_ppm1_n55);
   send_ppm1_sig_state_reg_2_inst : DF3 port map( D => send_ppm1_n95, C => 
                           i_clk_top, Q => send_ppm1_sig_state_2_port, QN => 
                           send_ppm1_n57);
   send_ppm1_sig_out_ppm_reg : DF3 port map( D => n132, C => i_clk_top, Q => 
                           o_ppm_top, QN => n_1000);
   send_ppm1_current_state_reg_2_inst : DF3 port map( D => n131, C => i_clk_top
                           , Q => send_ppm1_current_state_2_port, QN => n_1001)
                           ;
   send_ppm1_current_state_reg_1_inst : DF3 port map( D => send_ppm1_N82_port, 
                           C => i_clk_top, Q => send_ppm1_current_state_1_port,
                           QN => send_ppm1_n53);
   send_ppm1_sig_state_reg_0_inst : JK3 port map( J => send_ppm1_n69, K => n130
                           , C => i_clk_top, Q => send_ppm1_sig_state_0_port, 
                           QN => send_ppm1_n59);
   send_ppm1_local_counter1_o_count_reg_0_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N46, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_0_port, QN => n1);
   send_ppm1_local_counter1_o_count_reg_1_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N47, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_1_port, QN => n3);
   send_ppm1_local_counter1_o_count_reg_2_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N48, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_2_port, QN => n_1002);
   send_ppm1_local_counter1_o_count_reg_3_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N49, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_3_port, QN => n_1003);
   send_ppm1_local_counter1_o_count_reg_4_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N50, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_4_port, QN => n_1004);
   send_ppm1_local_counter1_o_count_reg_5_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N51, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_5_port, QN => n_1005);
   send_ppm1_local_counter1_o_count_reg_6_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N52, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_6_port, QN => n_1006);
   send_ppm1_local_counter1_o_count_reg_7_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N53, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_7_port, QN => n_1007);
   send_ppm1_local_counter1_o_count_reg_8_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N54, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_8_port, QN => n_1008);
   send_ppm1_local_counter1_o_count_reg_9_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N55, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_9_port, QN => n_1009);
   send_ppm1_local_counter1_o_count_reg_10_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N56, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_10_port, QN => n_1010)
                           ;
   send_ppm1_local_counter1_o_count_reg_11_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N57, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_11_port, QN => n_1011)
                           ;
   send_ppm1_local_counter1_o_count_reg_12_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N58, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_12_port, QN => n_1012)
                           ;
   send_ppm1_local_counter1_o_count_reg_13_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N59, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_13_port, QN => n_1013)
                           ;
   send_ppm1_local_counter1_o_count_reg_14_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N60, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_14_port, QN => n_1014)
                           ;
   send_ppm1_local_counter1_o_count_reg_15_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N61, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_15_port, QN => n_1015)
                           ;
   send_ppm1_local_counter1_o_count_reg_16_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N62, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_16_port, QN => n_1016)
                           ;
   send_ppm1_local_counter1_o_count_reg_17_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N63, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_17_port, QN => n_1017)
                           ;
   send_ppm1_local_counter1_o_count_reg_18_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N64, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_18_port, QN => n_1018)
                           ;
   send_ppm1_local_counter1_o_count_reg_19_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N65, C => i_clk_top, Q => 
                           send_ppm1_sig_out_local_count_19_port, QN => n_1019)
                           ;
   send_ppm1_local_counter1_v_val_reg_19_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N65, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_19_port, QN => n_1020
                           );
   send_ppm1_local_counter1_v_val_reg_18_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N64, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_18_port, QN => n_1021
                           );
   send_ppm1_local_counter1_v_val_reg_17_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N63, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_17_port, QN => n_1022
                           );
   send_ppm1_local_counter1_v_val_reg_16_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N62, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_16_port, QN => n_1023
                           );
   send_ppm1_local_counter1_v_val_reg_15_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N61, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_15_port, QN => n_1024
                           );
   send_ppm1_local_counter1_v_val_reg_14_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N60, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_14_port, QN => n_1025
                           );
   send_ppm1_local_counter1_v_val_reg_13_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N59, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_13_port, QN => n_1026
                           );
   send_ppm1_local_counter1_v_val_reg_12_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N58, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_12_port, QN => n_1027
                           );
   send_ppm1_local_counter1_v_val_reg_11_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N57, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_11_port, QN => n_1028
                           );
   send_ppm1_local_counter1_v_val_reg_10_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N56, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_10_port, QN => n_1029
                           );
   send_ppm1_local_counter1_v_val_reg_9_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N55, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_9_port, QN => n_1030)
                           ;
   send_ppm1_local_counter1_v_val_reg_8_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N54, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_8_port, QN => n_1031)
                           ;
   send_ppm1_local_counter1_v_val_reg_7_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N53, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_7_port, QN => n_1032)
                           ;
   send_ppm1_local_counter1_v_val_reg_6_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N52, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_6_port, QN => n_1033)
                           ;
   send_ppm1_local_counter1_v_val_reg_5_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N51, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_5_port, QN => n_1034)
                           ;
   send_ppm1_local_counter1_v_val_reg_4_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N50, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_4_port, QN => n_1035)
                           ;
   send_ppm1_local_counter1_v_val_reg_3_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N49, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_3_port, QN => n_1036)
                           ;
   send_ppm1_local_counter1_v_val_reg_2_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N48, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_2_port, QN => n_1037)
                           ;
   send_ppm1_local_counter1_v_val_reg_1_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N47, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_1_port, QN => n_1038)
                           ;
   send_ppm1_local_counter1_v_val_reg_0_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N46, C => i_clk_top, Q => 
                           send_ppm1_local_counter1_v_val_0_port, QN => n_1039)
                           ;
   send_ppm1_sig_reg_storage_reg_6_inst : DFE1 port map( D => n123, E => n127, 
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_6_port, QN => n_1040);
   send_ppm1_sig_reg_storage_reg_13_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n126, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_13_port, QN => n_1041);
   send_ppm1_sig_reg_storage_reg_14_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n126, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_14_port, QN => n_1042);
   send_ppm1_sig_reg_storage_reg_22_inst : DFE1 port map( D => n123, E => n125,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_22_port, QN => n_1043);
   send_ppm1_sig_reg_storage_reg_29_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n124, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_29_port, QN => n_1044);
   send_ppm1_sig_reg_storage_reg_30_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n124, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_30_port, QN => n_1045);
   send_ppm1_sig_reg_storage_reg_5_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n127, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_5_port, QN => n_1046);
   send_ppm1_sig_reg_storage_reg_21_inst : DFE1 port map( D => n123, E => n125,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_21_port, QN => n_1047);
   send_ppm1_sig_reg_storage_reg_12_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n126, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_12_port, QN => n8);
   send_ppm1_sig_reg_storage_reg_20_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n125, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_20_port, QN => n2);
   send_ppm1_sig_reg_storage_reg_28_inst : DFE1 port map( D => n123, E => n124,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_28_port, QN => n7);
   send_ppm1_sig_reg_storage_reg_3_inst : DFE1 port map( D => n123, E => n128, 
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_3_port, QN => n_1048);
   send_ppm1_sig_reg_storage_reg_10_inst : DFE1 port map( D => n123, E => n127,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_10_port, QN => n_1049);
   send_ppm1_sig_reg_storage_reg_11_inst : DFE1 port map( D => n123, E => n126,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_11_port, QN => n_1050);
   send_ppm1_sig_reg_storage_reg_18_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n125, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_18_port, QN => n_1051);
   send_ppm1_sig_reg_storage_reg_19_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n125, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_19_port, QN => n_1052);
   send_ppm1_sig_reg_storage_reg_26_inst : DFE1 port map( D => n123, E => n124,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_26_port, QN => n_1053);
   send_ppm1_sig_reg_storage_reg_27_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n124, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_27_port, QN => n_1054);
   send_ppm1_sig_reg_storage_reg_4_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n127, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_4_port, QN => n4);
   send_ppm1_sig_reg_storage_reg_2_inst : DFE1 port map( D => n123, E => n128, 
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_2_port, QN => n_1055);
   send_ppm1_sig_reg_storage_reg_23_inst : DFE1 port map( D => i_sel_top(1), E 
                           => n125, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_23_port, QN => n21);
   send_ppm1_sig_reg_storage_reg_15_inst : DFE1 port map( D => i_sel_top(1), E 
                           => n126, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_15_port, QN => n20);
   send_ppm1_sig_reg_storage_reg_31_inst : DFE1 port map( D => i_sel_top(1), E 
                           => n124, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_31_port, QN => n19);
   send_ppm1_sig_reg_storage_reg_7_inst : DFE1 port map( D => sig_reg_7_port, E
                           => n127, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_7_port, QN => n18);
   send_ppm1_sig_reg_storage_reg_9_inst : DFE1 port map( D => n123, E => n127, 
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_9_port, QN => n17);
   send_ppm1_sig_reg_storage_reg_17_inst : DFE1 port map( D => n123, E => n126,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_17_port, QN => n16);
   send_ppm1_sig_reg_storage_reg_25_inst : DFE1 port map( D => n123, E => n124,
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_25_port, QN => n15);
   send_ppm1_sig_reg_storage_reg_8_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n127, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_8_port, QN => n14);
   send_ppm1_sig_reg_storage_reg_16_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n126, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_16_port, QN => n13);
   send_ppm1_sig_reg_storage_reg_1_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n128, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_1_port, QN => n6);
   send_ppm1_sig_reg_storage_reg_24_inst : DFE1 port map( D => i_sel_top(0), E 
                           => n125, C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_24_port, QN => n22);
   send_ppm1_sig_reg_storage_reg_0_inst : DFE1 port map( D => n123, E => n128, 
                           C => i_clk_top, Q => 
                           send_ppm1_sig_reg_storage_0_port, QN => n9);
   U1 : NOR21 port map( A => n121, B => n24, Q => send_ppm1_local_counter1_N65)
                           ;
   U2 : MUX22 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, B 
                           => n150, S => 
                           send_ppm1_dp_cluster_1_mult_114_A2_8_port, Q => n5);
   U3 : MUX22 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, B 
                           => n192, S => 
                           send_ppm1_dp_cluster_4_mult_123_A2_8_port, Q => n10)
                           ;
   U4 : MUX22 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, B 
                           => n182, S => 
                           send_ppm1_dp_cluster_3_mult_120_A2_8_port, Q => n11)
                           ;
   U5 : MUX22 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, B 
                           => n170, S => 
                           send_ppm1_dp_cluster_2_mult_117_A2_8_port, Q => n12)
                           ;
   U6 : XNR21 port map( A => n143, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, Q 
                           => send_ppm1_dp_cluster_0_N279);
   U7 : XNR21 port map( A => send_ppm1_dp_cluster_0_N279, B => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, Q 
                           => send_ppm1_N196);
   U8 : INV3 port map( A => send_ppm1_dp_cluster_0_N48, Q => n166);
   U9 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, B 
                           => send_ppm1_dp_cluster_0_N279, Q => n55);
   U10 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_12_port, B => n60, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port);
   U11 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, Q 
                           => n60);
   U12 : INV3 port map( A => n53, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port);
   U13 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, B 
                           => n143, Q => n53);
   U14 : XNR21 port map( A => n143, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, Q 
                           => send_ppm1_dp_cluster_0_N280);
   U15 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_12_port, Q => n188);
   U16 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, B 
                           => n146, Q => send_ppm1_dp_cluster_0_N28);
   U17 : INV3 port map( A => send_ppm1_dp_cluster_0_N45, Q => n172);
   U18 : INV3 port map( A => send_ppm1_dp_cluster_0_N46, Q => n169);
   U19 : INV3 port map( A => send_ppm1_dp_cluster_0_N47, Q => n168);
   U20 : INV3 port map( A => send_ppm1_dp_cluster_0_N49, Q => n165);
   U21 : INV3 port map( A => n54, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port);
   U22 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, B 
                           => send_ppm1_dp_cluster_0_N280, Q => n54);
   U23 : INV3 port map( A => n52, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port);
   U24 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, B 
                           => n143, Q => n52);
   U25 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_13_port, B => n61, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port);
   U26 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, Q 
                           => n61);
   U27 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_11_port, B => n59, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port);
   U28 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, Q 
                           => n59);
   U29 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_10_port, B => n27, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port);
   U30 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_12_port, Q => n146);
   U31 : INV3 port map( A => n27, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port);
   U32 : NOR21 port map( A => n152, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, Q 
                           => n27);
   U33 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, Q 
                           => n143);
   U34 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, Q 
                           => n162);
   U35 : XNR21 port map( A => n143, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, Q 
                           => send_ppm1_dp_cluster_0_N281);
   U36 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_10_port, Q => n191);
   U37 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port, B 
                           => n149, Q => send_ppm1_dp_cluster_0_N26);
   U38 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_9_port, Q => n194);
   U39 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, B 
                           => n152, Q => send_ppm1_dp_cluster_0_N25);
   U40 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_13_port, Q => n187);
   U41 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, B 
                           => n145, Q => send_ppm1_dp_cluster_0_N29);
   U42 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_11_port, Q => n190);
   U43 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, B 
                           => n148, Q => send_ppm1_dp_cluster_0_N27);
   U44 : INV3 port map( A => send_ppm1_dp_cluster_0_N41, Q => n176);
   U45 : INV3 port map( A => send_ppm1_dp_cluster_0_N42, Q => n175);
   U46 : INV3 port map( A => send_ppm1_dp_cluster_0_N43, Q => n174);
   U47 : INV3 port map( A => send_ppm1_dp_cluster_0_N44, Q => n173);
   U48 : INV3 port map( A => send_ppm1_dp_cluster_0_N50, Q => n164);
   U49 : INV3 port map( A => send_ppm1_dp_cluster_0_N51, Q => n163);
   U50 : INV3 port map( A => n51, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port);
   U51 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, B 
                           => n143, Q => n51);
   U52 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_2_N250, Q => 
                           send_ppm1_sig_cyclesTrame2_12_port);
   U53 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_3_N235, Q => 
                           send_ppm1_sig_cyclesTrame3_12_port);
   U54 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_1_N265, Q => 
                           send_ppm1_sig_cyclesTrame1_12_port);
   U55 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_4_N220, Q => 
                           send_ppm1_sig_cyclesTrame4_12_port);
   U56 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_5_port, B => n58, Q =>
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port);
   U57 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, Q 
                           => n58);
   U58 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_8_port, B => n26, Q =>
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port);
   U59 : NOR21 port map( A => n102, B => n103, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port);
   U60 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, Q
                           => n102);
   U61 : INV3 port map( A => send_ppm1_dp_cluster_3_N235, Q => n103);
   U62 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_14_port, B => n62, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port);
   U63 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, Q 
                           => n62);
   U64 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_9_port, Q => n152);
   U65 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_13_port, Q => n145);
   U66 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_11_port, Q => n148);
   U67 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_10_port, Q => n149);
   U68 : NOR21 port map( A => n74, B => n75, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port);
   U69 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, Q
                           => n74);
   U70 : INV3 port map( A => send_ppm1_dp_cluster_1_N265, Q => n75);
   U71 : INV3 port map( A => n25, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port);
   U72 : NOR21 port map( A => n155, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, Q 
                           => n25);
   U73 : INV3 port map( A => n26, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port);
   U74 : NOR21 port map( A => n154, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, Q 
                           => n26);
   U75 : NOR21 port map( A => n88, B => n89, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port);
   U76 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, Q
                           => n88);
   U77 : INV3 port map( A => send_ppm1_dp_cluster_2_N250, Q => n89);
   U78 : NOR21 port map( A => n116, B => n117, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port);
   U79 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, Q
                           => n116);
   U80 : INV3 port map( A => send_ppm1_dp_cluster_4_N220, Q => n117);
   U81 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_15_port, B => n63, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port);
   U82 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, Q 
                           => n63);
   U83 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, B 
                           => n32, Q => send_ppm1_dp_cluster_0_N31);
   U84 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_6_port, Q => n197);
   U85 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, B 
                           => n155, Q => send_ppm1_dp_cluster_0_N22);
   U86 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_14_port, Q => n186);
   U87 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, B 
                           => n144, Q => send_ppm1_dp_cluster_0_N30);
   U88 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_5_port, Q => n198);
   U89 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, B 
                           => n156, Q => send_ppm1_dp_cluster_0_N21);
   U90 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_7_port, Q => n196);
   U91 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, B 
                           => n154, Q => send_ppm1_dp_cluster_0_N23);
   U92 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_8_port, Q => n195);
   U93 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port, B 
                           => n153, Q => send_ppm1_dp_cluster_0_N24);
   U94 : INV3 port map( A => send_ppm1_dp_cluster_0_N39, Q => n178);
   U95 : INV3 port map( A => send_ppm1_dp_cluster_0_N40, Q => n177);
   U96 : INV3 port map( A => send_ppm1_N198, Q => n141);
   U97 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port, 
                           B => send_ppm1_dp_cluster_2_N251, Q => 
                           send_ppm1_sig_cyclesTrame2_11_port);
   U98 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
                           B => send_ppm1_dp_cluster_3_N234, Q => 
                           send_ppm1_sig_cyclesTrame3_13_port);
   U99 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port, 
                           B => send_ppm1_dp_cluster_3_N236, Q => 
                           send_ppm1_sig_cyclesTrame3_11_port);
   U100 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_1_N268, Q => 
                           send_ppm1_sig_cyclesTrame1_9_port);
   U101 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port,
                           B => send_ppm1_dp_cluster_1_N264, Q => 
                           send_ppm1_sig_cyclesTrame1_13_port);
   U102 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port,
                           B => send_ppm1_dp_cluster_1_N266, Q => 
                           send_ppm1_sig_cyclesTrame1_11_port);
   U103 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port,
                           B => send_ppm1_dp_cluster_4_N221, Q => 
                           send_ppm1_sig_cyclesTrame4_11_port);
   U104 : XOR21 port map( A => n246, B => n147, Q => 
                           send_ppm1_dp_cluster_1_N265);
   U105 : XOR21 port map( A => n228, B => n189, Q => 
                           send_ppm1_dp_cluster_4_N220);
   U106 : XOR21 port map( A => n234, B => n181, Q => 
                           send_ppm1_dp_cluster_3_N235);
   U107 : XOR21 port map( A => n240, B => n167, Q => 
                           send_ppm1_dp_cluster_2_N250);
   U108 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port,
                           B => n5, Q => send_ppm1_sig_cyclesTrame1_10_port);
   U109 : NOR21 port map( A => n76, B => n77, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port);
   U110 : INV3 port map( A => send_ppm1_dp_cluster_1_N264, Q => n77);
   U111 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port, 
                           Q => n76);
   U112 : NOR21 port map( A => n46, B => n115, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port);
   U113 : INV3 port map( A => send_ppm1_dp_cluster_4_N221, Q => n115);
   U114 : NOR21 port map( A => n41, B => n101, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port);
   U115 : INV3 port map( A => send_ppm1_dp_cluster_3_N236, Q => n101);
   U116 : NOR21 port map( A => n36, B => n87, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port);
   U117 : INV3 port map( A => send_ppm1_dp_cluster_2_N251, Q => n87);
   U118 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_4_port, B => n57, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port);
   U119 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, Q 
                           => n57);
   U120 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_7_port, Q => n154);
   U121 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_8_port, Q => n153);
   U122 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_5_port, Q => n156);
   U123 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_6_port, Q => n155);
   U124 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_14_port, Q => n144);
   U125 : NOR21 port map( A => n71, B => n72, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port);
   U126 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, Q
                           => n71);
   U127 : INV3 port map( A => send_ppm1_dp_cluster_1_N268, Q => n72);
   U128 : NOR21 port map( A => n31, B => n73, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port);
   U129 : INV3 port map( A => send_ppm1_dp_cluster_1_N266, Q => n73);
   U130 : INV3 port map( A => n31, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port);
   U131 : NOR21 port map( A => n5, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port, Q 
                           => n31);
   U132 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port,
                           B => send_ppm1_dp_cluster_2_N249, Q => 
                           send_ppm1_sig_cyclesTrame2_13_port);
   U133 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_2_N253, Q => 
                           send_ppm1_sig_cyclesTrame2_9_port);
   U134 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_3_N238, Q => 
                           send_ppm1_sig_cyclesTrame3_9_port);
   U135 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port,
                           B => n12, Q => send_ppm1_sig_cyclesTrame2_10_port);
   U136 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port,
                           B => n11, Q => send_ppm1_sig_cyclesTrame3_10_port);
   U137 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port,
                           B => send_ppm1_dp_cluster_4_N219, Q => 
                           send_ppm1_sig_cyclesTrame4_13_port);
   U138 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_4_N223, Q => 
                           send_ppm1_sig_cyclesTrame4_9_port);
   U139 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port,
                           B => n10, Q => send_ppm1_sig_cyclesTrame4_10_port);
   U140 : NOR21 port map( A => n99, B => n100, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port);
   U141 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, Q
                           => n99);
   U142 : INV3 port map( A => send_ppm1_dp_cluster_3_N238, Q => n100);
   U143 : NOR21 port map( A => n85, B => n86, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port);
   U144 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, Q
                           => n85);
   U145 : INV3 port map( A => send_ppm1_dp_cluster_2_N253, Q => n86);
   U146 : NOR21 port map( A => n118, B => n119, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port);
   U147 : INV3 port map( A => send_ppm1_dp_cluster_4_N219, Q => n119);
   U148 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port, 
                           Q => n118);
   U149 : NOR21 port map( A => n104, B => n105, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port);
   U150 : INV3 port map( A => send_ppm1_dp_cluster_3_N234, Q => n105);
   U151 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
                           Q => n104);
   U152 : NOR21 port map( A => n90, B => n91, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port);
   U153 : INV3 port map( A => send_ppm1_dp_cluster_2_N249, Q => n91);
   U154 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port, 
                           Q => n90);
   U155 : INV3 port map( A => n46, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port);
   U156 : NOR21 port map( A => n10, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port, Q 
                           => n46);
   U157 : INV3 port map( A => n41, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port);
   U158 : NOR21 port map( A => n11, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port, Q 
                           => n41);
   U159 : INV3 port map( A => n36, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port);
   U160 : NOR21 port map( A => n12, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port, Q 
                           => n36);
   U161 : NOR21 port map( A => n113, B => n114, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port);
   U162 : INV3 port map( A => send_ppm1_dp_cluster_4_N223, Q => n114);
   U163 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, Q
                           => n113);
   U164 : BUF2 port map( A => n138, Q => n124);
   U165 : BUF2 port map( A => n138, Q => n125);
   U166 : BUF2 port map( A => n138, Q => n126);
   U167 : BUF2 port map( A => n138, Q => n127);
   U168 : BUF2 port map( A => n138, Q => n128);
   U169 : NOR40 port map( A => n142, B => n275, C => n274, D => n273, Q => 
                           send_ppm1_N198);
   U170 : NAND31 port map( A => n270, B => n269, C => n268, Q => n274);
   U171 : NAND22 port map( A => n272, B => n271, Q => n273);
   U172 : INV3 port map( A => n261, Q => n142);
   U173 : NAND41 port map( A => n161, B => n267, C => n266, D => n265, Q => 
                           n275);
   U174 : NAND22 port map( A => n3, B => send_ppm1_N179, Q => n267);
   U175 : INV3 port map( A => n262, Q => n161);
   U176 : NOR21 port map( A => n264, B => n263, Q => n265);
   U177 : NOR40 port map( A => n260, B => n259, C => n258, D => n257, Q => n261
                           );
   U178 : NAND31 port map( A => n249, B => n248, C => n247, Q => n260);
   U179 : NAND22 port map( A => n251, B => n250, Q => n259);
   U180 : NAND31 port map( A => n254, B => n253, C => n252, Q => n258);
   U181 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_3_port, B => n56, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port);
   U182 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, Q 
                           => n56);
   U183 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_3_port, Q => n200);
   U184 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, B 
                           => n158, Q => send_ppm1_dp_cluster_0_N19);
   U185 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_4_port, Q => n199);
   U186 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, B 
                           => n157, Q => send_ppm1_dp_cluster_0_N20);
   U187 : INV3 port map( A => n50, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port);
   U188 : INV3 port map( A => send_ppm1_dp_cluster_0_N38, Q => n179);
   U189 : NOR21 port map( A => n23, B => send_ppm1_dp_cluster_0_N296, Q => n50)
                           ;
   U190 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n121);
   U191 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n120);
   U192 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_2_port, Q => n159);
   U193 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_3_port, Q => n158);
   U194 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_4_port, Q => n157);
   U195 : NOR21 port map( A => n121, B => n206, Q => 
                           send_ppm1_local_counter1_N63);
   U196 : INV3 port map( A => send_ppm1_local_counter1_N23, Q => n206);
   U197 : NOR21 port map( A => n121, B => n208, Q => 
                           send_ppm1_local_counter1_N61);
   U198 : INV3 port map( A => send_ppm1_local_counter1_N21, Q => n208);
   U199 : NOR21 port map( A => n121, B => n210, Q => 
                           send_ppm1_local_counter1_N59);
   U200 : INV3 port map( A => send_ppm1_local_counter1_N19, Q => n210);
   U201 : NOR21 port map( A => n121, B => n212, Q => 
                           send_ppm1_local_counter1_N57);
   U202 : INV3 port map( A => send_ppm1_local_counter1_N17, Q => n212);
   U203 : NOR21 port map( A => n121, B => n214, Q => 
                           send_ppm1_local_counter1_N55);
   U204 : INV3 port map( A => send_ppm1_local_counter1_N15, Q => n214);
   U205 : NOR21 port map( A => n121, B => n216, Q => 
                           send_ppm1_local_counter1_N53);
   U206 : INV3 port map( A => send_ppm1_local_counter1_N13, Q => n216);
   U207 : NOR21 port map( A => n120, B => n217, Q => 
                           send_ppm1_local_counter1_N52);
   U208 : INV3 port map( A => send_ppm1_local_counter1_N12, Q => n217);
   U209 : NOR21 port map( A => n120, B => n218, Q => 
                           send_ppm1_local_counter1_N51);
   U210 : INV3 port map( A => send_ppm1_local_counter1_N11, Q => n218);
   U211 : NOR21 port map( A => n120, B => n219, Q => 
                           send_ppm1_local_counter1_N50);
   U212 : INV3 port map( A => send_ppm1_local_counter1_N10, Q => n219);
   U213 : NOR21 port map( A => n120, B => n220, Q => 
                           send_ppm1_local_counter1_N49);
   U214 : INV3 port map( A => send_ppm1_local_counter1_N9, Q => n220);
   U215 : NOR21 port map( A => n120, B => n221, Q => 
                           send_ppm1_local_counter1_N48);
   U216 : INV3 port map( A => send_ppm1_local_counter1_N8, Q => n221);
   U217 : NOR21 port map( A => n120, B => n222, Q => 
                           send_ppm1_local_counter1_N47);
   U218 : INV3 port map( A => send_ppm1_local_counter1_N7, Q => n222);
   U219 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_5_port);
   U220 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_8_port);
   U221 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_5_port);
   U222 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_8_port);
   U223 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_8_port);
   U224 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_5_port);
   U225 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_5_port);
   U226 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_7_port);
   U227 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_7_port);
   U228 : XOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_A1_11_port, B =>
                           n245, Q => send_ppm1_dp_cluster_1_N264);
   U229 : NOR21 port map( A => n147, B => n246, Q => n245);
   U230 : XOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_1_N268);
   U231 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_1_N263, Q => 
                           send_ppm1_sig_cyclesTrame1_14_port);
   U232 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_6_port);
   U233 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_6_port);
   U234 : XOR21 port map( A => n151, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_1_N266);
   U235 : XOR21 port map( A => n193, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_4_N221);
   U236 : XOR21 port map( A => n183, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_3_N236);
   U237 : XOR21 port map( A => n171, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_2_N251);
   U238 : NAND22 port map( A => n151, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           n246);
   U239 : NOR21 port map( A => n29, B => n67, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port);
   U240 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, Q 
                           => n67);
   U241 : NOR21 port map( A => n64, B => n65, Q => 
                           send_ppm1_dp_cluster_1_mult_114_A2_8_port);
   U242 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, Q 
                           => n65);
   U243 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           Q => n64);
   U244 : NOR21 port map( A => n69, B => n70, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port);
   U245 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, Q
                           => n69);
   U246 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, Q 
                           => n70);
   U247 : NOR21 port map( A => n30, B => n68, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port);
   U248 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, Q 
                           => n68);
   U249 : INV3 port map( A => n49, Q => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port);
   U250 : NOR21 port map( A => n13, B => n14, Q => n49);
   U251 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port, Q 
                           => n147);
   U252 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port, Q 
                           => n189);
   U253 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port, Q 
                           => n181);
   U254 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port, Q 
                           => n167);
   U255 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, Q 
                           => n150);
   U256 : INV3 port map( A => n241, Q => n151);
   U257 : NAND22 port map( A => send_ppm1_dp_cluster_1_mult_114_A2_8_port, B =>
                           send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, Q => 
                           n241);
   U258 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n122);
   U259 : XOR21 port map( A => n14, B => n13, Q => n23);
   U260 : INV3 port map( A => n30, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port);
   U261 : NOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, Q
                           => n30);
   U262 : NOR21 port map( A => n122, B => n205, Q => 
                           send_ppm1_local_counter1_N64);
   U263 : INV3 port map( A => send_ppm1_local_counter1_N24, Q => n205);
   U264 : NOR21 port map( A => n122, B => n207, Q => 
                           send_ppm1_local_counter1_N62);
   U265 : INV3 port map( A => send_ppm1_local_counter1_N22_port, Q => n207);
   U266 : NOR21 port map( A => n122, B => n209, Q => 
                           send_ppm1_local_counter1_N60);
   U267 : INV3 port map( A => send_ppm1_local_counter1_N20, Q => n209);
   U268 : NOR21 port map( A => n122, B => n211, Q => 
                           send_ppm1_local_counter1_N58);
   U269 : INV3 port map( A => send_ppm1_local_counter1_N18, Q => n211);
   U270 : NOR21 port map( A => n122, B => n213, Q => 
                           send_ppm1_local_counter1_N56);
   U271 : INV3 port map( A => send_ppm1_local_counter1_N16, Q => n213);
   U272 : NOR21 port map( A => n122, B => n215, Q => 
                           send_ppm1_local_counter1_N54);
   U273 : INV3 port map( A => send_ppm1_local_counter1_N14, Q => n215);
   U274 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_8_port);
   U275 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_7_port);
   U276 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_7_port);
   U277 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_2_N248, Q => 
                           send_ppm1_sig_cyclesTrame2_14_port);
   U278 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_6_port);
   U279 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_3_N233, Q => 
                           send_ppm1_sig_cyclesTrame3_14_port);
   U280 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_6_port);
   U281 : XOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_A1_11_port, B =>
                           n227, Q => send_ppm1_dp_cluster_4_N219);
   U282 : NOR21 port map( A => n189, B => n228, Q => n227);
   U283 : XOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_A1_11_port, B =>
                           n233, Q => send_ppm1_dp_cluster_3_N234);
   U284 : NOR21 port map( A => n181, B => n234, Q => n233);
   U285 : XOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_A1_11_port, B =>
                           n239, Q => send_ppm1_dp_cluster_2_N249);
   U286 : NOR21 port map( A => n167, B => n240, Q => n239);
   U287 : XOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_4_N223);
   U288 : XOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_3_N238);
   U289 : XOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_2_N253);
   U290 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_4_N218, Q => 
                           send_ppm1_sig_cyclesTrame4_14_port);
   U291 : NAND22 port map( A => n193, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           n228);
   U292 : NAND22 port map( A => n183, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           n234);
   U293 : NAND22 port map( A => n171, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           n240);
   U294 : NOR21 port map( A => n44, B => n109, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port);
   U295 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, Q 
                           => n109);
   U296 : NOR21 port map( A => n39, B => n95, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port);
   U297 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, Q 
                           => n95);
   U298 : NOR21 port map( A => n34, B => n81, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port);
   U299 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, Q 
                           => n81);
   U300 : NOR21 port map( A => n106, B => n107, Q => 
                           send_ppm1_dp_cluster_4_mult_123_A2_8_port);
   U301 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, Q 
                           => n107);
   U302 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           Q => n106);
   U303 : NOR21 port map( A => n111, B => n112, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port);
   U304 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, Q
                           => n111);
   U305 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, Q 
                           => n112);
   U306 : NOR21 port map( A => n97, B => n98, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port);
   U307 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, Q
                           => n97);
   U308 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, Q 
                           => n98);
   U309 : NOR21 port map( A => n83, B => n84, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port);
   U310 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, Q
                           => n83);
   U311 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, Q 
                           => n84);
   U312 : NOR21 port map( A => n45, B => n110, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port);
   U313 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, Q 
                           => n110);
   U314 : NOR21 port map( A => n40, B => n96, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port);
   U315 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, Q 
                           => n96);
   U316 : NOR21 port map( A => n35, B => n82, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port);
   U317 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, Q 
                           => n82);
   U318 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, Q 
                           => n192);
   U319 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, Q 
                           => n182);
   U320 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, Q 
                           => n170);
   U321 : INV3 port map( A => n223, Q => n193);
   U322 : NAND22 port map( A => send_ppm1_dp_cluster_4_mult_123_A2_8_port, B =>
                           send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, Q => 
                           n223);
   U323 : INV3 port map( A => n229, Q => n183);
   U324 : NAND22 port map( A => send_ppm1_dp_cluster_3_mult_120_A2_8_port, B =>
                           send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, Q => 
                           n229);
   U325 : INV3 port map( A => n235, Q => n171);
   U326 : NAND22 port map( A => send_ppm1_dp_cluster_2_mult_117_A2_8_port, B =>
                           send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, Q => 
                           n235);
   U327 : NOR21 port map( A => n147, B => n244, Q => n243);
   U328 : NAND22 port map( A => n151, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           n244);
   U329 : NOR21 port map( A => n189, B => n226, Q => n225);
   U330 : NAND22 port map( A => n193, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           n226);
   U331 : NOR21 port map( A => n181, B => n232, Q => n231);
   U332 : NAND22 port map( A => n183, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           n232);
   U333 : NOR21 port map( A => n167, B => n238, Q => n237);
   U334 : NAND22 port map( A => n171, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           n238);
   U335 : INV3 port map( A => n32, Q => send_ppm1_sig_cyclesTrame1_15_port);
   U336 : NOR21 port map( A => send_ppm1_dp_cluster_1_N263, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port, Q 
                           => n32);
   U337 : INV3 port map( A => n45, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port);
   U338 : NOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, Q
                           => n45);
   U339 : INV3 port map( A => n40, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port);
   U340 : NOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, Q
                           => n40);
   U341 : INV3 port map( A => n35, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port);
   U342 : NOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, Q
                           => n35);
   U343 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, 
                           Q => n66);
   U344 : NOR21 port map( A => n92, B => n93, Q => 
                           send_ppm1_dp_cluster_3_mult_120_A2_8_port);
   U345 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           Q => n92);
   U346 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, Q 
                           => n93);
   U347 : NOR21 port map( A => n78, B => n79, Q => 
                           send_ppm1_dp_cluster_2_mult_117_A2_8_port);
   U348 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           Q => n78);
   U349 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, Q 
                           => n79);
   U350 : INV3 port map( A => n37, Q => send_ppm1_sig_cyclesTrame2_15_port);
   U351 : NOR21 port map( A => send_ppm1_dp_cluster_2_N248, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port, Q 
                           => n37);
   U352 : INV3 port map( A => n42, Q => send_ppm1_sig_cyclesTrame3_15_port);
   U353 : NOR21 port map( A => send_ppm1_dp_cluster_3_N233, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port, Q 
                           => n42);
   U354 : INV3 port map( A => n47, Q => send_ppm1_sig_cyclesTrame4_15_port);
   U355 : NOR21 port map( A => send_ppm1_dp_cluster_4_N218, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port, Q 
                           => n47);
   U356 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, 
                           Q => n108);
   U357 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, 
                           Q => n94);
   U358 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, 
                           Q => n80);
   U359 : NOR40 port map( A => n363, B => n362, C => n361, D => n360, Q => 
                           send_ppm1_N148);
   U360 : NAND41 port map( A => n160, B => n347, C => n346, D => n345, Q => 
                           n363);
   U361 : NAND41 port map( A => n351, B => n350, C => n349, D => n348, Q => 
                           n362);
   U362 : NAND41 port map( A => n355, B => n354, C => n353, D => n352, Q => 
                           n361);
   U363 : XNR21 port map( A => send_ppm1_dp_cluster_0_N296, B => n23, Q => 
                           send_ppm1_N179);
   U364 : AOI221 port map( A => n3, B => n1, C => n1, D => send_ppm1_N179, Q =>
                           n262);
   U365 : NOR21 port map( A => n3, B => n13, Q => n298);
   U366 : NOR21 port map( A => n3, B => n14, Q => n320);
   U367 : INV3 port map( A => n342, Q => n160);
   U368 : NOR21 port map( A => n3, B => n9, Q => n342);
   U369 : NOR21 port map( A => n3, B => n22, Q => n276);
   U370 : NOR31 port map( A => send_ppm1_n71, B => send_ppm1_n72, C => 
                           send_ppm1_n70, Q => send_ppm1_n69);
   U371 : INV3 port map( A => send_ppm1_n71, Q => n203);
   U372 : INV3 port map( A => send_ppm1_n72, Q => n137);
   U373 : INV3 port map( A => send_ppm1_n76, Q => n140);
   U374 : INV3 port map( A => send_ppm1_n60, Q => n138);
   U375 : INV3 port map( A => send_ppm1_n70, Q => n132);
   U376 : BUF2 port map( A => sig_reg_28_port, Q => n123);
   U377 : NOR21 port map( A => n135, B => n134, Q => sig_reg_28_port);
   U378 : NAND22 port map( A => n135, B => n134, Q => sig_reg_7_port);
   U379 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => 
                           send_ppm1_sig_reg_storage_1_port, Q => 
                           send_ppm1_sig_cyclesTrame1_2_port);
   U380 : INV3 port map( A => send_ppm1_n73, Q => n130);
   U381 : OAI2111 port map( A => n203, B => send_ppm1_n70, C => send_ppm1_n74, 
                           D => send_ppm1_n75, Q => send_ppm1_n73);
   U382 : NAND31 port map( A => send_ppm1_n63, B => send_ppm1_n53, C => 
                           i_reset_n_top, Q => send_ppm1_n75);
   U383 : NAND31 port map( A => send_ppm1_n76, B => n141, C => i_reset_n_top, Q
                           => send_ppm1_n74);
   U384 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_2_port, Q => 
                           send_ppm1_sig_cyclesTrame1_3_port);
   U385 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_3_port, Q => 
                           send_ppm1_sig_cyclesTrame1_4_port);
   U386 : NAND22 port map( A => send_ppm1_sig_state_0_port, B => send_ppm1_n58,
                           Q => send_ppm1_n65);
   U387 : INV3 port map( A => send_ppm1_n69, Q => n133);
   U388 : INV3 port map( A => send_ppm1_n66, Q => n129);
   U389 : NOR21 port map( A => n9, B => n6, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port);
   U390 : NOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, B
                           => n9, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port);
   U391 : NAND41 port map( A => send_ppm1_n69, B => send_ppm1_sig_state_1_port,
                           C => send_ppm1_sig_state_0_port, D => send_ppm1_n57,
                           Q => send_ppm1_n68);
   U392 : AOI211 port map( A => n132, B => send_ppm1_n58, C => send_ppm1_n66, Q
                           => send_ppm1_n67);
   U393 : XNR21 port map( A => send_ppm1_N194, B => 
                           send_ppm1_sig_out_local_count_16_port, Q => n252);
   U394 : INV3 port map( A => n48, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port);
   U395 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_2_port, Q => n201);
   U396 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => n159, Q 
                           => send_ppm1_dp_cluster_0_N18);
   U397 : NAND22 port map( A => i_reset_n_top, B => n136, Q => 
                           send_ppm1_local_counter1_n22);
   U398 : INV3 port map( A => send_ppm1_sig_in_init, Q => n136);
   U399 : OAI2111 port map( A => n140, B => n141, C => send_ppm1_n60, D => 
                           send_ppm1_n61, Q => send_ppm1_sig_in_init);
   U400 : AOI221 port map( A => n203, B => send_ppm1_n62, C => send_ppm1_n63, D
                           => send_ppm1_n64, Q => send_ppm1_n61);
   U401 : XNR21 port map( A => send_ppm1_N197, B => 
                           send_ppm1_sig_out_local_count_19_port, Q => n266);
   U402 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port, B 
                           => send_ppm1_dp_cluster_0_N278, Q => send_ppm1_N197)
                           ;
   U403 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port, B 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, Q 
                           => send_ppm1_dp_cluster_0_N278);
   U404 : INV3 port map( A => n55, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port);
   U405 : INV3 port map( A => n28, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port);
   U406 : NOR21 port map( A => send_ppm1_sig_reg_storage_2_port, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, Q =>
                           n28);
   U407 : NAND22 port map( A => n256, B => n255, Q => n257);
   U408 : XNR21 port map( A => send_ppm1_N195, B => 
                           send_ppm1_sig_out_local_count_17_port, Q => n255);
   U409 : XNR21 port map( A => send_ppm1_N196, B => 
                           send_ppm1_sig_out_local_count_18_port, Q => n256);
   U410 : XNR21 port map( A => send_ppm1_dp_cluster_0_N280, B => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, Q 
                           => send_ppm1_N195);
   U411 : NOR21 port map( A => n120, B => send_ppm1_local_counter1_v_val_0_port
                           , Q => send_ppm1_local_counter1_N46);
   U412 : XNR21 port map( A => send_ppm1_local_counter1_add_34_carry_19_port, B
                           => send_ppm1_local_counter1_v_val_19_port, Q => n24)
                           ;
   U413 : XOR21 port map( A => send_ppm1_sig_reg_storage_8_port, B => 
                           send_ppm1_sig_reg_storage_9_port, Q => 
                           send_ppm1_sig_cyclesTrame2_2_port);
   U414 : XOR21 port map( A => send_ppm1_sig_reg_storage_16_port, B => 
                           send_ppm1_sig_reg_storage_17_port, Q => 
                           send_ppm1_sig_cyclesTrame3_2_port);
   U415 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_10_port, Q => 
                           send_ppm1_sig_cyclesTrame2_3_port);
   U416 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_11_port, Q => 
                           send_ppm1_sig_cyclesTrame2_4_port);
   U417 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_18_port, Q => 
                           send_ppm1_sig_cyclesTrame3_3_port);
   U418 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_19_port, Q => 
                           send_ppm1_sig_cyclesTrame3_4_port);
   U419 : XOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => 
                           send_ppm1_sig_reg_storage_25_port, Q => 
                           send_ppm1_sig_cyclesTrame4_2_port);
   U420 : XOR21 port map( A => send_ppm1_sig_reg_storage_4_port, B => 
                           send_ppm1_sig_reg_storage_0_port, Q => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port);
   U421 : XNR21 port map( A => n242, B => 
                           send_ppm1_dp_cluster_1_mult_114_A2_12_port, Q => 
                           send_ppm1_dp_cluster_1_N263);
   U422 : NOR21 port map( A => n66, B => n18, Q => 
                           send_ppm1_dp_cluster_1_mult_114_A2_12_port);
   U423 : NAND22 port map( A => send_ppm1_dp_cluster_1_mult_114_A1_11_port, B 
                           => n243, Q => n242);
   U424 : XNR21 port map( A => n9, B => send_ppm1_sig_reg_storage_24_port, Q =>
                           send_ppm1_dp_cluster_0_N296);
   U425 : XOR21 port map( A => send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_1_mult_114_A1_11_port);
   U426 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_26_port, Q => 
                           send_ppm1_sig_cyclesTrame4_3_port);
   U427 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_27_port, Q => 
                           send_ppm1_sig_cyclesTrame4_4_port);
   U428 : NOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => n9, Q =>
                           n48);
   U429 : NOR21 port map( A => n22, B => n15, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port);
   U430 : NOR21 port map( A => n22, B => n15, Q => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port);
   U431 : NOR21 port map( A => n9, B => n6, Q => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port);
   U432 : NOR21 port map( A => n7, B => n22, Q => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port);
   U433 : XOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => 
                           send_ppm1_sig_reg_storage_25_port, Q => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port);
   U434 : NOR21 port map( A => n4, B => n9, Q => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port);
   U435 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => 
                           send_ppm1_sig_reg_storage_1_port, Q => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port);
   U436 : NOR21 port map( A => n13, B => n16, Q => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port);
   U437 : NOR21 port map( A => n14, B => n17, Q => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port);
   U438 : NOR21 port map( A => n2, B => n13, Q => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port);
   U439 : XOR21 port map( A => send_ppm1_sig_reg_storage_16_port, B => 
                           send_ppm1_sig_reg_storage_17_port, Q => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port);
   U440 : NOR21 port map( A => n13, B => n16, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port);
   U441 : NOR21 port map( A => n14, B => n17, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port);
   U442 : XNR21 port map( A => send_ppm1_N193, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n254);
   U443 : INV3 port map( A => n43, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port);
   U444 : NOR21 port map( A => send_ppm1_sig_reg_storage_26_port, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, Q =>
                           n43);
   U445 : INV3 port map( A => n38, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port);
   U446 : NOR21 port map( A => send_ppm1_sig_reg_storage_18_port, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, Q =>
                           n38);
   U447 : INV3 port map( A => n33, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port);
   U448 : NOR21 port map( A => send_ppm1_sig_reg_storage_10_port, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, Q =>
                           n33);
   U449 : INV3 port map( A => n29, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port);
   U450 : NOR21 port map( A => send_ppm1_sig_reg_storage_3_port, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, Q =>
                           n29);
   U451 : INV3 port map( A => n44, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port);
   U452 : NOR21 port map( A => send_ppm1_sig_reg_storage_27_port, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, Q =>
                           n44);
   U453 : INV3 port map( A => n39, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port);
   U454 : NOR21 port map( A => send_ppm1_sig_reg_storage_19_port, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, Q =>
                           n39);
   U455 : INV3 port map( A => n34, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port);
   U456 : NOR21 port map( A => send_ppm1_sig_reg_storage_11_port, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, Q =>
                           n34);
   U457 : INV3 port map( A => send_ppm1_n77, Q => n131);
   U458 : NAND31 port map( A => i_reset_n_top, B => send_ppm1_n76, C => 
                           send_ppm1_N198, Q => send_ppm1_n77);
   U459 : XOR21 port map( A => send_ppm1_sig_reg_storage_28_port, B => 
                           send_ppm1_sig_reg_storage_24_port, Q => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port);
   U460 : XOR21 port map( A => send_ppm1_sig_reg_storage_20_port, B => 
                           send_ppm1_sig_reg_storage_16_port, Q => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port);
   U461 : XOR21 port map( A => send_ppm1_sig_reg_storage_12_port, B => 
                           send_ppm1_sig_reg_storage_8_port, Q => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port);
   U462 : XNR21 port map( A => n224, B => 
                           send_ppm1_dp_cluster_4_mult_123_A2_12_port, Q => 
                           send_ppm1_dp_cluster_4_N218);
   U463 : NOR21 port map( A => n108, B => n19, Q => 
                           send_ppm1_dp_cluster_4_mult_123_A2_12_port);
   U464 : NAND22 port map( A => send_ppm1_dp_cluster_4_mult_123_A1_11_port, B 
                           => n225, Q => n224);
   U465 : XNR21 port map( A => n236, B => 
                           send_ppm1_dp_cluster_2_mult_117_A2_12_port, Q => 
                           send_ppm1_dp_cluster_2_N248);
   U466 : NOR21 port map( A => n80, B => n20, Q => 
                           send_ppm1_dp_cluster_2_mult_117_A2_12_port);
   U467 : NAND22 port map( A => send_ppm1_dp_cluster_2_mult_117_A1_11_port, B 
                           => n237, Q => n236);
   U468 : XOR21 port map( A => send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_4_mult_123_A1_11_port);
   U469 : XOR21 port map( A => send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_3_mult_120_A1_11_port);
   U470 : XOR21 port map( A => send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_2_mult_117_A1_11_port);
   U471 : OAI2111 port map( A => send_ppm1_N198, B => n140, C => send_ppm1_n78,
                           D => i_reset_n_top, Q => send_ppm1_N82_port);
   U472 : NAND31 port map( A => send_ppm1_n72, B => n203, C => send_ppm1_n79, Q
                           => send_ppm1_n78);
   U473 : NOR21 port map( A => n8, B => n14, Q => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port);
   U474 : XOR21 port map( A => send_ppm1_sig_reg_storage_8_port, B => 
                           send_ppm1_sig_reg_storage_9_port, Q => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port);
   U475 : XNR21 port map( A => send_ppm1_N192, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n253);
   U476 : XNR21 port map( A => n230, B => 
                           send_ppm1_dp_cluster_3_mult_120_A2_12_port, Q => 
                           send_ppm1_dp_cluster_3_N233);
   U477 : NOR21 port map( A => n94, B => n21, Q => 
                           send_ppm1_dp_cluster_3_mult_120_A2_12_port);
   U478 : NAND22 port map( A => send_ppm1_dp_cluster_3_mult_120_A1_11_port, B 
                           => n231, Q => n230);
   U479 : XNR21 port map( A => send_ppm1_N190, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n250);
   U480 : XNR21 port map( A => send_ppm1_N191, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n251);
   U481 : XNR21 port map( A => send_ppm1_N189, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n247);
   U482 : XNR21 port map( A => send_ppm1_N188, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n249);
   U483 : XNR21 port map( A => send_ppm1_N187, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n248);
   U484 : NAND41 port map( A => n334, B => n337, C => n336, D => n335, Q => 
                           n338);
   U485 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n334);
   U486 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n335);
   U487 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n337);
   U488 : NAND41 port map( A => n312, B => n315, C => n314, D => n313, Q => 
                           n316);
   U489 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n312);
   U490 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n313);
   U491 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n315);
   U492 : NAND41 port map( A => n356, B => n359, C => n358, D => n357, Q => 
                           n360);
   U493 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n356);
   U494 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n357);
   U495 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n359);
   U496 : INV3 port map( A => send_ppm1_N169, Q => n185);
   U497 : AOI311 port map( A => send_ppm1_N148, B => send_ppm1_n58, C => 
                           send_ppm1_sig_state_0_port, D => send_ppm1_n92, Q =>
                           send_ppm1_n91);
   U498 : NOR40 port map( A => n297, B => n296, C => n295, D => n294, Q => 
                           send_ppm1_N169);
   U499 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n336);
   U500 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n314);
   U501 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n358);
   U502 : NOR21 port map( A => send_ppm1_n93, B => send_ppm1_n58, Q => 
                           send_ppm1_n92);
   U503 : AOI221 port map( A => send_ppm1_N156, B => send_ppm1_n59, C => 
                           send_ppm1_N163, D => send_ppm1_sig_state_0_port, Q 
                           => send_ppm1_n93);
   U504 : NOR40 port map( A => n319, B => n318, C => n317, D => n316, Q => 
                           send_ppm1_N163);
   U505 : NOR40 port map( A => n341, B => n340, C => n339, D => n338, Q => 
                           send_ppm1_N156);
   U506 : NAND41 port map( A => n290, B => n293, C => n292, D => n291, Q => 
                           n294);
   U507 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n290);
   U508 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n291);
   U509 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n293);
   U510 : NAND41 port map( A => n333, B => n332, C => n331, D => n330, Q => 
                           n339);
   U511 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n330);
   U512 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n331);
   U513 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n332);
   U514 : NAND41 port map( A => n311, B => n310, C => n309, D => n308, Q => 
                           n317);
   U515 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n308);
   U516 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n309);
   U517 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n310);
   U518 : NAND41 port map( A => n289, B => n288, C => n287, D => n286, Q => 
                           n295);
   U519 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n286);
   U520 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n287);
   U521 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n288);
   U522 : OAI2111 port map( A => send_ppm1_n64, B => send_ppm1_n80, C => 
                           send_ppm1_n81, D => i_reset_n_top, Q => 
                           send_ppm1_N81_port);
   U523 : NAND22 port map( A => send_ppm1_n63, B => send_ppm1_n53, Q => 
                           send_ppm1_n80);
   U524 : NAND31 port map( A => n203, B => n137, C => send_ppm1_n79, Q => 
                           send_ppm1_n81);
   U525 : XNR21 port map( A => send_ppm1_N185, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n271);
   U526 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n333);
   U527 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n311);
   U528 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n355);
   U529 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n289);
   U530 : XNR21 port map( A => send_ppm1_N186, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n272);
   U531 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n292);
   U532 : XNR21 port map( A => send_ppm1_N184, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n268);
   U533 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n354);
   U534 : NAND41 port map( A => n329, B => n328, C => n327, D => n326, Q => 
                           n340);
   U535 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n326);
   U536 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n327);
   U537 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n328);
   U538 : NAND41 port map( A => n307, B => n306, C => n305, D => n304, Q => 
                           n318);
   U539 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n304);
   U540 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n305);
   U541 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n306);
   U542 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n329);
   U543 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n307);
   U544 : XNR21 port map( A => send_ppm1_N182, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n269);
   U545 : XNR21 port map( A => send_ppm1_N183, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n270);
   U546 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n353);
   U547 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n352);
   U548 : NAND41 port map( A => n285, B => n284, C => n283, D => n282, Q => 
                           n296);
   U549 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n282);
   U550 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n283);
   U551 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n284);
   U552 : XOR21 port map( A => send_ppm1_N180, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n264);
   U553 : XOR21 port map( A => send_ppm1_N181, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n263);
   U554 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n351);
   U555 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n285);
   U556 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n350);
   U557 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n349);
   U558 : NAND41 port map( A => n180, B => n325, C => n324, D => n323, Q => 
                           n341);
   U559 : INV3 port map( A => n320, Q => n180);
   U560 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n324);
   U561 : NAND41 port map( A => n184, B => n303, C => n302, D => n301, Q => 
                           n319);
   U562 : INV3 port map( A => n298, Q => n184);
   U563 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n302);
   U564 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n348);
   U565 : NOR21 port map( A => n322, B => n321, Q => n323);
   U566 : XOR21 port map( A => send_ppm1_sig_cyclesTrame2_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n322);
   U567 : XOR21 port map( A => send_ppm1_sig_cyclesTrame2_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n321);
   U568 : NOR21 port map( A => n300, B => n299, Q => n301);
   U569 : XOR21 port map( A => send_ppm1_sig_cyclesTrame3_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n300);
   U570 : XOR21 port map( A => send_ppm1_sig_cyclesTrame3_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n299);
   U571 : NOR21 port map( A => n344, B => n343, Q => n345);
   U572 : XOR21 port map( A => send_ppm1_sig_cyclesTrame1_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n344);
   U573 : XOR21 port map( A => send_ppm1_sig_cyclesTrame1_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n343);
   U574 : NAND41 port map( A => n202, B => n281, C => n280, D => n279, Q => 
                           n297);
   U575 : INV3 port map( A => n276, Q => n202);
   U576 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n280);
   U577 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n346);
   U578 : NOR21 port map( A => n278, B => n277, Q => n279);
   U579 : XOR21 port map( A => send_ppm1_sig_cyclesTrame4_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n278);
   U580 : XOR21 port map( A => send_ppm1_sig_cyclesTrame4_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n277);
   U581 : NAND41 port map( A => send_ppm1_n82, B => send_ppm1_n83, C => 
                           send_ppm1_n84, D => send_ppm1_n85, Q => 
                           send_ppm1_n71);
   U582 : NOR21 port map( A => send_ppm1_sig_out_local_count_16_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => 
                           send_ppm1_n82);
   U583 : NOR31 port map( A => send_ppm1_sig_out_local_count_17_port, B => 
                           send_ppm1_sig_out_local_count_19_port, C => 
                           send_ppm1_sig_out_local_count_18_port, Q => 
                           send_ppm1_n83);
   U584 : NOR40 port map( A => send_ppm1_sig_out_local_count_5_port, B => n204,
                           C => send_ppm1_sig_out_local_count_4_port, D => 
                           send_ppm1_sig_out_local_count_2_port, Q => 
                           send_ppm1_n84);
   U585 : NOR31 port map( A => send_ppm1_sig_state_0_port, B => 
                           send_ppm1_sig_state_1_port, C => send_ppm1_n57, Q =>
                           send_ppm1_n72);
   U586 : NOR31 port map( A => send_ppm1_n86, B => send_ppm1_n87, C => 
                           send_ppm1_n88, Q => send_ppm1_n85);
   U587 : NAND22 port map( A => send_ppm1_sig_out_local_count_8_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => 
                           send_ppm1_n88);
   U588 : NAND31 port map( A => send_ppm1_sig_out_local_count_1_port, B => 
                           send_ppm1_sig_out_local_count_12_port, C => 
                           send_ppm1_sig_out_local_count_3_port, Q => 
                           send_ppm1_n87);
   U589 : NAND41 port map( A => send_ppm1_sig_out_local_count_11_port, B => 
                           send_ppm1_sig_out_local_count_10_port, C => 
                           send_ppm1_n89, D => 
                           send_ppm1_sig_out_local_count_0_port, Q => 
                           send_ppm1_n86);
   U590 : NOR21 port map( A => send_ppm1_sig_out_local_count_14_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => 
                           send_ppm1_n89);
   U591 : INV3 port map( A => send_ppm1_n90, Q => n204);
   U592 : NOR21 port map( A => send_ppm1_sig_out_local_count_9_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => 
                           send_ppm1_n90);
   U593 : NOR31 port map( A => send_ppm1_current_state_0_port, B => 
                           send_ppm1_current_state_2_port, C => send_ppm1_n53, 
                           Q => send_ppm1_n76);
   U594 : AOI221 port map( A => send_ppm1_n63, B => 
                           send_ppm1_current_state_1_port, C => send_ppm1_n62, 
                           D => send_ppm1_current_state_2_port, Q => 
                           send_ppm1_n60);
   U595 : NAND22 port map( A => i_reset_n_top, B => send_ppm1_n79, Q => 
                           send_ppm1_n70);
   U596 : NOR21 port map( A => send_ppm1_n55, B => 
                           send_ppm1_current_state_2_port, Q => send_ppm1_n63);
   U597 : NOR21 port map( A => send_ppm1_current_state_0_port, B => 
                           send_ppm1_current_state_1_port, Q => send_ppm1_n62);
   U598 : NOR21 port map( A => n139, B => send_ppm1_current_state_2_port, Q => 
                           send_ppm1_n79);
   U599 : INV3 port map( A => send_ppm1_n62, Q => n139);
   U600 : INV3 port map( A => i_sel_top(1), Q => n134);
   U601 : INV3 port map( A => i_sel_top(0), Q => n135);
   U602 : OAI222 port map( A => n1, B => n3, C => n22, D => n1, Q => n281);
   U603 : OAI222 port map( A => n1, B => n3, C => n13, D => n1, Q => n303);
   U604 : OAI222 port map( A => n1, B => n3, C => n14, D => n1, Q => n325);
   U605 : OAI222 port map( A => n1, B => n3, C => n9, D => n1, Q => n347);

end SYN_rtl;
