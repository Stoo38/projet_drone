
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_top_ppm is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_top_ppm;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_top_ppm.all;

entity top_ppm is

   port( i_clk_top, i_reset_n_top : in std_logic;  i_sel_top : in 
         std_logic_vector (3 downto 0);  o_ppm_top : out std_logic);

end top_ppm;

architecture SYN_rtl of top_ppm is

   component OAI222
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component BUF2
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component INV3
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component XNR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI2111
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR21
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR40
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI221
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND22
      port( A, B : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND41
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI211
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI311
      port( A, B, C, D : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR31
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   component BUF6
      port( A : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX22
      port( A, B, S : in std_logic;  Q : out std_logic);
   end component;
   
   component DFE1
      port( D, E, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DF3
      port( D, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component JK3
      port( J, K, C : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component ADD32
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADD22
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI212
      port( A, B, C : in std_logic;  Q : out std_logic);
   end component;
   
   signal sig_clk25, N3, sig_reg_31_port, sig_reg_30_port, sig_reg_22_port, 
      sig_reg_15_port, sig_reg_14_port, sig_reg_7_port, sig_reg_6_port, 
      decoder1_n14, decoder1_n13, decoder1_n12, decoder1_n11, decoder1_n10, 
      decoder1_n9, decoder1_n8, send_ppm1_n95, send_ppm1_n94, send_ppm1_n93, 
      send_ppm1_n92, send_ppm1_n91, send_ppm1_n90, send_ppm1_n89, send_ppm1_n88
      , send_ppm1_n87, send_ppm1_n86, send_ppm1_n85, send_ppm1_n84, 
      send_ppm1_n83, send_ppm1_n82, send_ppm1_n81, send_ppm1_n80, send_ppm1_n79
      , send_ppm1_n78, send_ppm1_n77, send_ppm1_n76, send_ppm1_n75, 
      send_ppm1_n74, send_ppm1_n73, send_ppm1_n72, send_ppm1_n71, send_ppm1_n70
      , send_ppm1_n69, send_ppm1_n68, send_ppm1_n67, send_ppm1_n66, 
      send_ppm1_n65, send_ppm1_n64, send_ppm1_n63, send_ppm1_n62, send_ppm1_n61
      , send_ppm1_n60, send_ppm1_n59, send_ppm1_n58, send_ppm1_n57, 
      send_ppm1_n55, send_ppm1_n53, send_ppm1_dp_cluster_4_N218, 
      send_ppm1_dp_cluster_4_N219, send_ppm1_dp_cluster_4_N220, 
      send_ppm1_dp_cluster_4_N221, send_ppm1_dp_cluster_4_N223, 
      send_ppm1_dp_cluster_3_N233, send_ppm1_dp_cluster_3_N234, 
      send_ppm1_dp_cluster_3_N235, send_ppm1_dp_cluster_3_N236, 
      send_ppm1_dp_cluster_3_N238, send_ppm1_dp_cluster_2_N248, 
      send_ppm1_dp_cluster_2_N249, send_ppm1_dp_cluster_2_N250, 
      send_ppm1_dp_cluster_2_N251, send_ppm1_dp_cluster_2_N253, 
      send_ppm1_dp_cluster_1_N263, send_ppm1_dp_cluster_1_N264, 
      send_ppm1_dp_cluster_1_N265, send_ppm1_dp_cluster_1_N266, 
      send_ppm1_dp_cluster_1_N268, send_ppm1_dp_cluster_0_N18, 
      send_ppm1_dp_cluster_0_N19, send_ppm1_dp_cluster_0_N20, 
      send_ppm1_dp_cluster_0_N21, send_ppm1_dp_cluster_0_N22, 
      send_ppm1_dp_cluster_0_N23, send_ppm1_dp_cluster_0_N24, 
      send_ppm1_dp_cluster_0_N25, send_ppm1_dp_cluster_0_N26, 
      send_ppm1_dp_cluster_0_N27, send_ppm1_dp_cluster_0_N278, 
      send_ppm1_dp_cluster_0_N279, send_ppm1_dp_cluster_0_N28, 
      send_ppm1_dp_cluster_0_N280, send_ppm1_dp_cluster_0_N281, 
      send_ppm1_dp_cluster_0_N282, send_ppm1_dp_cluster_0_N283, 
      send_ppm1_dp_cluster_0_N284, send_ppm1_dp_cluster_0_N285, 
      send_ppm1_dp_cluster_0_N286, send_ppm1_dp_cluster_0_N287, 
      send_ppm1_dp_cluster_0_N288, send_ppm1_dp_cluster_0_N289, 
      send_ppm1_dp_cluster_0_N29, send_ppm1_dp_cluster_0_N290, 
      send_ppm1_dp_cluster_0_N291, send_ppm1_dp_cluster_0_N292, 
      send_ppm1_dp_cluster_0_N293, send_ppm1_dp_cluster_0_N294, 
      send_ppm1_dp_cluster_0_N295, send_ppm1_dp_cluster_0_N296, 
      send_ppm1_dp_cluster_0_N30, send_ppm1_dp_cluster_0_N31, 
      send_ppm1_dp_cluster_0_N38, send_ppm1_dp_cluster_0_N39, 
      send_ppm1_dp_cluster_0_N40, send_ppm1_dp_cluster_0_N41, 
      send_ppm1_dp_cluster_0_N42, send_ppm1_dp_cluster_0_N43, 
      send_ppm1_dp_cluster_0_N44, send_ppm1_dp_cluster_0_N45, 
      send_ppm1_dp_cluster_0_N46, send_ppm1_dp_cluster_0_N47, 
      send_ppm1_dp_cluster_0_N48, send_ppm1_dp_cluster_0_N49, 
      send_ppm1_dp_cluster_0_N50, send_ppm1_dp_cluster_0_N51, send_ppm1_N198, 
      send_ppm1_N197, send_ppm1_N196, send_ppm1_N195, send_ppm1_N194, 
      send_ppm1_N193, send_ppm1_N192, send_ppm1_N191, send_ppm1_N190, 
      send_ppm1_N189, send_ppm1_N188, send_ppm1_N187, send_ppm1_N186, 
      send_ppm1_N185, send_ppm1_N184, send_ppm1_N183, send_ppm1_N182, 
      send_ppm1_N181, send_ppm1_N180, send_ppm1_N179, send_ppm1_N169, 
      send_ppm1_N163, send_ppm1_N156, send_ppm1_N148, send_ppm1_N82_port, 
      send_ppm1_N81_port, send_ppm1_sig_state_0_port, 
      send_ppm1_sig_state_1_port, send_ppm1_sig_state_2_port, 
      send_ppm1_current_state_0_port, send_ppm1_current_state_1_port, 
      send_ppm1_current_state_2_port, send_ppm1_sig_cyclesTrame4_2_port, 
      send_ppm1_sig_cyclesTrame4_3_port, send_ppm1_sig_cyclesTrame4_4_port, 
      send_ppm1_sig_cyclesTrame4_5_port, send_ppm1_sig_cyclesTrame4_6_port, 
      send_ppm1_sig_cyclesTrame4_7_port, send_ppm1_sig_cyclesTrame4_8_port, 
      send_ppm1_sig_cyclesTrame4_9_port, send_ppm1_sig_cyclesTrame4_10_port, 
      send_ppm1_sig_cyclesTrame4_11_port, send_ppm1_sig_cyclesTrame4_12_port, 
      send_ppm1_sig_cyclesTrame4_13_port, send_ppm1_sig_cyclesTrame4_14_port, 
      send_ppm1_sig_cyclesTrame4_15_port, send_ppm1_sig_cyclesTrame3_2_port, 
      send_ppm1_sig_cyclesTrame3_3_port, send_ppm1_sig_cyclesTrame3_4_port, 
      send_ppm1_sig_cyclesTrame3_5_port, send_ppm1_sig_cyclesTrame3_6_port, 
      send_ppm1_sig_cyclesTrame3_7_port, send_ppm1_sig_cyclesTrame3_8_port, 
      send_ppm1_sig_cyclesTrame3_9_port, send_ppm1_sig_cyclesTrame3_10_port, 
      send_ppm1_sig_cyclesTrame3_11_port, send_ppm1_sig_cyclesTrame3_12_port, 
      send_ppm1_sig_cyclesTrame3_13_port, send_ppm1_sig_cyclesTrame3_14_port, 
      send_ppm1_sig_cyclesTrame3_15_port, send_ppm1_sig_cyclesTrame2_2_port, 
      send_ppm1_sig_cyclesTrame2_3_port, send_ppm1_sig_cyclesTrame2_4_port, 
      send_ppm1_sig_cyclesTrame2_5_port, send_ppm1_sig_cyclesTrame2_6_port, 
      send_ppm1_sig_cyclesTrame2_7_port, send_ppm1_sig_cyclesTrame2_8_port, 
      send_ppm1_sig_cyclesTrame2_9_port, send_ppm1_sig_cyclesTrame2_10_port, 
      send_ppm1_sig_cyclesTrame2_11_port, send_ppm1_sig_cyclesTrame2_12_port, 
      send_ppm1_sig_cyclesTrame2_13_port, send_ppm1_sig_cyclesTrame2_14_port, 
      send_ppm1_sig_cyclesTrame2_15_port, send_ppm1_sig_cyclesTrame1_2_port, 
      send_ppm1_sig_cyclesTrame1_3_port, send_ppm1_sig_cyclesTrame1_4_port, 
      send_ppm1_sig_cyclesTrame1_5_port, send_ppm1_sig_cyclesTrame1_6_port, 
      send_ppm1_sig_cyclesTrame1_7_port, send_ppm1_sig_cyclesTrame1_8_port, 
      send_ppm1_sig_cyclesTrame1_9_port, send_ppm1_sig_cyclesTrame1_10_port, 
      send_ppm1_sig_cyclesTrame1_11_port, send_ppm1_sig_cyclesTrame1_12_port, 
      send_ppm1_sig_cyclesTrame1_13_port, send_ppm1_sig_cyclesTrame1_14_port, 
      send_ppm1_sig_cyclesTrame1_15_port, send_ppm1_sig_reg_storage_0_port, 
      send_ppm1_sig_reg_storage_1_port, send_ppm1_sig_reg_storage_2_port, 
      send_ppm1_sig_reg_storage_3_port, send_ppm1_sig_reg_storage_4_port, 
      send_ppm1_sig_reg_storage_5_port, send_ppm1_sig_reg_storage_6_port, 
      send_ppm1_sig_reg_storage_7_port, send_ppm1_sig_reg_storage_8_port, 
      send_ppm1_sig_reg_storage_9_port, send_ppm1_sig_reg_storage_10_port, 
      send_ppm1_sig_reg_storage_11_port, send_ppm1_sig_reg_storage_12_port, 
      send_ppm1_sig_reg_storage_13_port, send_ppm1_sig_reg_storage_14_port, 
      send_ppm1_sig_reg_storage_15_port, send_ppm1_sig_reg_storage_16_port, 
      send_ppm1_sig_reg_storage_17_port, send_ppm1_sig_reg_storage_18_port, 
      send_ppm1_sig_reg_storage_19_port, send_ppm1_sig_reg_storage_20_port, 
      send_ppm1_sig_reg_storage_21_port, send_ppm1_sig_reg_storage_22_port, 
      send_ppm1_sig_reg_storage_23_port, send_ppm1_sig_reg_storage_24_port, 
      send_ppm1_sig_reg_storage_25_port, send_ppm1_sig_reg_storage_26_port, 
      send_ppm1_sig_reg_storage_27_port, send_ppm1_sig_reg_storage_28_port, 
      send_ppm1_sig_reg_storage_29_port, send_ppm1_sig_reg_storage_30_port, 
      send_ppm1_sig_reg_storage_31_port, send_ppm1_sig_out_local_count_0_port, 
      send_ppm1_sig_out_local_count_1_port, 
      send_ppm1_sig_out_local_count_2_port, 
      send_ppm1_sig_out_local_count_3_port, 
      send_ppm1_sig_out_local_count_4_port, 
      send_ppm1_sig_out_local_count_5_port, 
      send_ppm1_sig_out_local_count_6_port, 
      send_ppm1_sig_out_local_count_7_port, 
      send_ppm1_sig_out_local_count_8_port, 
      send_ppm1_sig_out_local_count_9_port, 
      send_ppm1_sig_out_local_count_10_port, 
      send_ppm1_sig_out_local_count_11_port, 
      send_ppm1_sig_out_local_count_12_port, 
      send_ppm1_sig_out_local_count_13_port, 
      send_ppm1_sig_out_local_count_14_port, 
      send_ppm1_sig_out_local_count_15_port, 
      send_ppm1_sig_out_local_count_16_port, 
      send_ppm1_sig_out_local_count_17_port, 
      send_ppm1_sig_out_local_count_18_port, 
      send_ppm1_sig_out_local_count_19_port, send_ppm1_sig_in_init, 
      send_ppm1_local_counter1_n22, send_ppm1_local_counter1_N65, 
      send_ppm1_local_counter1_N64, send_ppm1_local_counter1_N63, 
      send_ppm1_local_counter1_N62, send_ppm1_local_counter1_N61, 
      send_ppm1_local_counter1_N60, send_ppm1_local_counter1_N59, 
      send_ppm1_local_counter1_N58, send_ppm1_local_counter1_N57, 
      send_ppm1_local_counter1_N56, send_ppm1_local_counter1_N55, 
      send_ppm1_local_counter1_N54, send_ppm1_local_counter1_N53, 
      send_ppm1_local_counter1_N52, send_ppm1_local_counter1_N51, 
      send_ppm1_local_counter1_N50, send_ppm1_local_counter1_N49, 
      send_ppm1_local_counter1_N48, send_ppm1_local_counter1_N47, 
      send_ppm1_local_counter1_N46, send_ppm1_local_counter1_N24, 
      send_ppm1_local_counter1_N23, send_ppm1_local_counter1_N22_port, 
      send_ppm1_local_counter1_N21, send_ppm1_local_counter1_N20, 
      send_ppm1_local_counter1_N19, send_ppm1_local_counter1_N18, 
      send_ppm1_local_counter1_N17, send_ppm1_local_counter1_N16, 
      send_ppm1_local_counter1_N15, send_ppm1_local_counter1_N14, 
      send_ppm1_local_counter1_N13, send_ppm1_local_counter1_N12, 
      send_ppm1_local_counter1_N11, send_ppm1_local_counter1_N10, 
      send_ppm1_local_counter1_N9, send_ppm1_local_counter1_N8, 
      send_ppm1_local_counter1_N7, send_ppm1_local_counter1_v_val_0_port, 
      send_ppm1_local_counter1_v_val_1_port, 
      send_ppm1_local_counter1_v_val_2_port, 
      send_ppm1_local_counter1_v_val_3_port, 
      send_ppm1_local_counter1_v_val_4_port, 
      send_ppm1_local_counter1_v_val_5_port, 
      send_ppm1_local_counter1_v_val_6_port, 
      send_ppm1_local_counter1_v_val_7_port, 
      send_ppm1_local_counter1_v_val_8_port, 
      send_ppm1_local_counter1_v_val_9_port, 
      send_ppm1_local_counter1_v_val_10_port, 
      send_ppm1_local_counter1_v_val_11_port, 
      send_ppm1_local_counter1_v_val_12_port, 
      send_ppm1_local_counter1_v_val_13_port, 
      send_ppm1_local_counter1_v_val_14_port, 
      send_ppm1_local_counter1_v_val_15_port, 
      send_ppm1_local_counter1_v_val_16_port, 
      send_ppm1_local_counter1_v_val_17_port, 
      send_ppm1_local_counter1_v_val_18_port, 
      send_ppm1_local_counter1_v_val_19_port, 
      send_ppm1_local_counter1_add_34_carry_2_port, 
      send_ppm1_local_counter1_add_34_carry_3_port, 
      send_ppm1_local_counter1_add_34_carry_4_port, 
      send_ppm1_local_counter1_add_34_carry_5_port, 
      send_ppm1_local_counter1_add_34_carry_6_port, 
      send_ppm1_local_counter1_add_34_carry_7_port, 
      send_ppm1_local_counter1_add_34_carry_8_port, 
      send_ppm1_local_counter1_add_34_carry_9_port, 
      send_ppm1_local_counter1_add_34_carry_10_port, 
      send_ppm1_local_counter1_add_34_carry_11_port, 
      send_ppm1_local_counter1_add_34_carry_12_port, 
      send_ppm1_local_counter1_add_34_carry_13_port, 
      send_ppm1_local_counter1_add_34_carry_14_port, 
      send_ppm1_local_counter1_add_34_carry_15_port, 
      send_ppm1_local_counter1_add_34_carry_16_port, 
      send_ppm1_local_counter1_add_34_carry_17_port, 
      send_ppm1_local_counter1_add_34_carry_18_port, 
      send_ppm1_local_counter1_add_34_carry_19_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, 
      send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, 
      send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port, 
      send_ppm1_dp_cluster_1_mult_114_A2_8_port, 
      send_ppm1_dp_cluster_1_mult_114_A2_12_port, 
      send_ppm1_dp_cluster_1_mult_114_A1_11_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, 
      send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port, 
      send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port, 
      send_ppm1_dp_cluster_2_mult_117_A2_8_port, 
      send_ppm1_dp_cluster_2_mult_117_A2_12_port, 
      send_ppm1_dp_cluster_2_mult_117_A1_11_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, 
      send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port, 
      send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port, 
      send_ppm1_dp_cluster_3_mult_120_A2_8_port, 
      send_ppm1_dp_cluster_3_mult_120_A2_12_port, 
      send_ppm1_dp_cluster_3_mult_120_A1_11_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, 
      send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
      send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port, 
      send_ppm1_dp_cluster_4_mult_123_A2_8_port, 
      send_ppm1_dp_cluster_4_mult_123_A2_12_port, 
      send_ppm1_dp_cluster_4_mult_123_A1_11_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, 
      send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
      send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port, 
      send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port, n2, n3_port, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, 
      n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, 
      n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, 
      n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, 
      n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, 
      n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056 : std_logic;

begin
   
   send_ppm1_U39 : OAI222 port map( A => n145, B => n193, C => 
                           send_ppm1_sig_state_2_port, D => send_ppm1_n91, Q =>
                           send_ppm1_n64);
   send_ppm1_U16 : OAI212 port map( A => send_ppm1_sig_state_0_port, B => 
                           send_ppm1_n70, C => n133, Q => send_ppm1_n66);
   send_ppm1_U13 : OAI212 port map( A => send_ppm1_n67, B => send_ppm1_n57, C 
                           => send_ppm1_n68, Q => send_ppm1_n95);
   send_ppm1_U6 : OAI222 port map( A => n132, B => send_ppm1_n58, C => n136, D 
                           => send_ppm1_n65, Q => send_ppm1_n94);
   send_ppm1_local_counter1_add_34_U1_1_1 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_1_port, B => 
                           send_ppm1_local_counter1_v_val_0_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_2_port, S => 
                           send_ppm1_local_counter1_N7);
   send_ppm1_local_counter1_add_34_U1_1_2 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_2_port, B => 
                           send_ppm1_local_counter1_add_34_carry_2_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_3_port, S => 
                           send_ppm1_local_counter1_N8);
   send_ppm1_local_counter1_add_34_U1_1_3 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_3_port, B => 
                           send_ppm1_local_counter1_add_34_carry_3_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_4_port, S => 
                           send_ppm1_local_counter1_N9);
   send_ppm1_local_counter1_add_34_U1_1_4 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_4_port, B => 
                           send_ppm1_local_counter1_add_34_carry_4_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_5_port, S => 
                           send_ppm1_local_counter1_N10);
   send_ppm1_local_counter1_add_34_U1_1_5 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_5_port, B => 
                           send_ppm1_local_counter1_add_34_carry_5_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_6_port, S => 
                           send_ppm1_local_counter1_N11);
   send_ppm1_local_counter1_add_34_U1_1_6 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_6_port, B => 
                           send_ppm1_local_counter1_add_34_carry_6_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_7_port, S => 
                           send_ppm1_local_counter1_N12);
   send_ppm1_local_counter1_add_34_U1_1_7 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_7_port, B => 
                           send_ppm1_local_counter1_add_34_carry_7_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_8_port, S => 
                           send_ppm1_local_counter1_N13);
   send_ppm1_local_counter1_add_34_U1_1_8 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_8_port, B => 
                           send_ppm1_local_counter1_add_34_carry_8_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_9_port, S => 
                           send_ppm1_local_counter1_N14);
   send_ppm1_local_counter1_add_34_U1_1_9 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_9_port, B => 
                           send_ppm1_local_counter1_add_34_carry_9_port, CO => 
                           send_ppm1_local_counter1_add_34_carry_10_port, S => 
                           send_ppm1_local_counter1_N15);
   send_ppm1_local_counter1_add_34_U1_1_10 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_10_port, B => 
                           send_ppm1_local_counter1_add_34_carry_10_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_11_port, S => 
                           send_ppm1_local_counter1_N16);
   send_ppm1_local_counter1_add_34_U1_1_11 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_11_port, B => 
                           send_ppm1_local_counter1_add_34_carry_11_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_12_port, S => 
                           send_ppm1_local_counter1_N17);
   send_ppm1_local_counter1_add_34_U1_1_12 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_12_port, B => 
                           send_ppm1_local_counter1_add_34_carry_12_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_13_port, S => 
                           send_ppm1_local_counter1_N18);
   send_ppm1_local_counter1_add_34_U1_1_13 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_13_port, B => 
                           send_ppm1_local_counter1_add_34_carry_13_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_14_port, S => 
                           send_ppm1_local_counter1_N19);
   send_ppm1_local_counter1_add_34_U1_1_14 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_14_port, B => 
                           send_ppm1_local_counter1_add_34_carry_14_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_15_port, S => 
                           send_ppm1_local_counter1_N20);
   send_ppm1_local_counter1_add_34_U1_1_15 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_15_port, B => 
                           send_ppm1_local_counter1_add_34_carry_15_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_16_port, S => 
                           send_ppm1_local_counter1_N21);
   send_ppm1_local_counter1_add_34_U1_1_16 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_16_port, B => 
                           send_ppm1_local_counter1_add_34_carry_16_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_17_port, S => 
                           send_ppm1_local_counter1_N22_port);
   send_ppm1_local_counter1_add_34_U1_1_17 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_17_port, B => 
                           send_ppm1_local_counter1_add_34_carry_17_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_18_port, S => 
                           send_ppm1_local_counter1_N23);
   send_ppm1_local_counter1_add_34_U1_1_18 : ADD22 port map( A => 
                           send_ppm1_local_counter1_v_val_18_port, B => 
                           send_ppm1_local_counter1_add_34_carry_18_port, CO =>
                           send_ppm1_local_counter1_add_34_carry_19_port, S => 
                           send_ppm1_local_counter1_N24);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_2 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_2_port, B => 
                           send_ppm1_sig_cyclesTrame3_2_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_dp_cluster_0_N38);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_3 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_3_port, B => 
                           send_ppm1_sig_cyclesTrame3_3_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_dp_cluster_0_N39);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_4 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_4_port, B => 
                           send_ppm1_sig_cyclesTrame3_4_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_dp_cluster_0_N40);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_5 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_5_port, B => 
                           send_ppm1_sig_cyclesTrame3_5_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_dp_cluster_0_N41);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_6 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_6_port, B => 
                           send_ppm1_sig_cyclesTrame3_6_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_dp_cluster_0_N42);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_7 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_7_port, B => 
                           send_ppm1_sig_cyclesTrame3_7_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_dp_cluster_0_N43);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_8 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_8_port, B => 
                           send_ppm1_sig_cyclesTrame3_8_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_dp_cluster_0_N44);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_9 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_9_port, B => 
                           send_ppm1_sig_cyclesTrame3_9_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_dp_cluster_0_N45);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_10 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_10_port, B => 
                           send_ppm1_sig_cyclesTrame3_10_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_dp_cluster_0_N46);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_11 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_11_port, B => 
                           send_ppm1_sig_cyclesTrame3_11_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_dp_cluster_0_N47);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_12 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_12_port, B => 
                           send_ppm1_sig_cyclesTrame3_12_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_dp_cluster_0_N48);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_13 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_13_port, B => 
                           send_ppm1_sig_cyclesTrame3_13_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_dp_cluster_0_N49);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_14 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_14_port, B => 
                           send_ppm1_sig_cyclesTrame3_14_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_dp_cluster_0_N50);
   send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_U1_15 : ADD32 port map( A => 
                           send_ppm1_sig_cyclesTrame2_15_port, B => 
                           send_ppm1_sig_cyclesTrame3_15_port, CI => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_dp_cluster_0_N51);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_2 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N18, B => n209, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_dp_cluster_0_N295);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_3 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N19, B => n208, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_dp_cluster_0_N294);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_4 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N20, B => n207, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_dp_cluster_0_N293);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_5 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N21, B => n206, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_dp_cluster_0_N292);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_6 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N22, B => n205, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_dp_cluster_0_N291);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_7 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N23, B => n204, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_dp_cluster_0_N290);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_8 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N24, B => n203, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_dp_cluster_0_N289);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_9 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N25, B => n202, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_dp_cluster_0_N288);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_10 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N26, B => n199, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_dp_cluster_0_N287);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_11 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N27, B => n198, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_dp_cluster_0_N286);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_12 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N28, B => n196, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_dp_cluster_0_N285);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_13 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N29, B => n195, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_dp_cluster_0_N284);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_14 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N30, B => n194, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_dp_cluster_0_N283);
   send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_U1_15 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N31, B => n48, CI => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_dp_cluster_0_N282);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_2 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N295, B => n187, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, S 
                           => send_ppm1_N180);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_3 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N294, B => n186, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_3_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, S 
                           => send_ppm1_N181);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_4 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N293, B => n185, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_4_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, S 
                           => send_ppm1_N182);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_5 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N292, B => n184, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_5_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, S 
                           => send_ppm1_N183);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_6 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N291, B => n183, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_6_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, S 
                           => send_ppm1_N184);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_7 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N290, B => n182, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_7_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, S 
                           => send_ppm1_N185);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_8 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N289, B => n181, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_8_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, S 
                           => send_ppm1_N186);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_9 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N288, B => n180, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_9_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, S 
                           => send_ppm1_N187);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_10 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N287, B => n177, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_10_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, S 
                           => send_ppm1_N188);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_11 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N286, B => n176, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_11_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, S 
                           => send_ppm1_N189);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_12 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N285, B => n174, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_12_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, S 
                           => send_ppm1_N190);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_13 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N284, B => n173, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_13_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, S 
                           => send_ppm1_N191);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_14 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N283, B => n172, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_14_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, S 
                           => send_ppm1_N192);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_15 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N282, B => n171, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_15_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, S 
                           => send_ppm1_N193);
   send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_U2_16 : ADD32 port map( A => 
                           send_ppm1_dp_cluster_0_N281, B => n170, CI => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_16_port, 
                           CO => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, S 
                           => send_ppm1_N194);
   send_ppm1_dp_cluster_1_mult_114_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_2_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_1_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_3_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_2_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_4_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_3_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port);
   send_ppm1_dp_cluster_1_mult_114_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_5_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_4_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port);
   send_ppm1_dp_cluster_1_mult_114_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_5_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port);
   send_ppm1_dp_cluster_1_mult_114_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_6_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_5_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port);
   send_ppm1_dp_cluster_1_mult_114_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_6_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port);
   send_ppm1_dp_cluster_1_mult_114_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_6_port, CO => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port);
   send_ppm1_dp_cluster_1_mult_114_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_1_mult_114_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port);
   send_ppm1_dp_cluster_2_mult_117_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_10_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_9_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_11_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_10_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_12_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_11_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port);
   send_ppm1_dp_cluster_2_mult_117_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_13_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_12_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port);
   send_ppm1_dp_cluster_2_mult_117_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_13_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port);
   send_ppm1_dp_cluster_2_mult_117_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_14_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_13_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port);
   send_ppm1_dp_cluster_2_mult_117_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_14_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port);
   send_ppm1_dp_cluster_2_mult_117_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_14_port, CO => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port);
   send_ppm1_dp_cluster_2_mult_117_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_2_mult_117_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port);
   send_ppm1_dp_cluster_3_mult_120_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_18_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_17_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_19_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_18_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_20_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_19_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port);
   send_ppm1_dp_cluster_3_mult_120_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_21_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_20_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port);
   send_ppm1_dp_cluster_3_mult_120_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_21_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port);
   send_ppm1_dp_cluster_3_mult_120_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_22_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_21_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port);
   send_ppm1_dp_cluster_3_mult_120_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_22_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port);
   send_ppm1_dp_cluster_3_mult_120_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_22_port, CO => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port);
   send_ppm1_dp_cluster_3_mult_120_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_3_mult_120_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port);
   send_ppm1_dp_cluster_4_mult_123_S3_2_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_26_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port, CI 
                           => send_ppm1_sig_reg_storage_25_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_3_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_27_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_2_5_port, CI 
                           => send_ppm1_sig_reg_storage_26_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_4_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_28_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_3_5_port, CI 
                           => send_ppm1_sig_reg_storage_27_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port);
   send_ppm1_dp_cluster_4_mult_123_S3_5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_29_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_5_port, CI 
                           => send_ppm1_sig_reg_storage_28_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port);
   send_ppm1_dp_cluster_4_mult_123_S2_5_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_29_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port);
   send_ppm1_dp_cluster_4_mult_123_S3_6_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_30_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_5_port, CI 
                           => send_ppm1_sig_reg_storage_29_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port);
   send_ppm1_dp_cluster_4_mult_123_S2_6_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_30_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_5_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_2_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port);
   send_ppm1_dp_cluster_4_mult_123_S5_5 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_5_port, CI 
                           => send_ppm1_sig_reg_storage_30_port, CO => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, S 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port);
   send_ppm1_dp_cluster_4_mult_123_S4_1 : ADD32 port map( A => 
                           send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_6_1_port, CI 
                           => send_ppm1_dp_cluster_4_mult_123_SUMB_3_5_port, CO
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           S => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port);
   sig_clk25_reg : DF3 port map( D => N3, C => i_clk_top, Q => sig_clk25, QN =>
                           n_1000);
   send_ppm1_sig_state_reg_1_inst : DF3 port map( D => send_ppm1_n94, C => n129
                           , Q => send_ppm1_sig_state_1_port, QN => 
                           send_ppm1_n58);
   send_ppm1_current_state_reg_0_inst : DF3 port map( D => send_ppm1_N81_port, 
                           C => n130, Q => send_ppm1_current_state_0_port, QN 
                           => send_ppm1_n55);
   send_ppm1_sig_state_reg_2_inst : DF3 port map( D => send_ppm1_n95, C => n130
                           , Q => send_ppm1_sig_state_2_port, QN => 
                           send_ppm1_n57);
   send_ppm1_sig_out_ppm_reg : DF3 port map( D => n135, C => n130, Q => 
                           o_ppm_top, QN => n_1001);
   send_ppm1_current_state_reg_2_inst : DF3 port map( D => n134, C => n130, Q 
                           => send_ppm1_current_state_2_port, QN => n_1002);
   send_ppm1_current_state_reg_1_inst : DF3 port map( D => send_ppm1_N82_port, 
                           C => n130, Q => send_ppm1_current_state_1_port, QN 
                           => send_ppm1_n53);
   send_ppm1_sig_state_reg_0_inst : JK3 port map( J => send_ppm1_n69, K => n133
                           , C => sig_clk25, Q => send_ppm1_sig_state_0_port, 
                           QN => send_ppm1_n59);
   send_ppm1_local_counter1_o_count_reg_0_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N46, C => n130, Q => 
                           send_ppm1_sig_out_local_count_0_port, QN => n3_port)
                           ;
   send_ppm1_local_counter1_o_count_reg_1_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N47, C => n130, Q => 
                           send_ppm1_sig_out_local_count_1_port, QN => n7);
   send_ppm1_local_counter1_o_count_reg_2_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N48, C => n130, Q => 
                           send_ppm1_sig_out_local_count_2_port, QN => n_1003);
   send_ppm1_local_counter1_o_count_reg_3_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N49, C => n130, Q => 
                           send_ppm1_sig_out_local_count_3_port, QN => n_1004);
   send_ppm1_local_counter1_o_count_reg_4_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N50, C => n130, Q => 
                           send_ppm1_sig_out_local_count_4_port, QN => n_1005);
   send_ppm1_local_counter1_o_count_reg_5_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N51, C => n129, Q => 
                           send_ppm1_sig_out_local_count_5_port, QN => n_1006);
   send_ppm1_local_counter1_o_count_reg_6_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N52, C => n129, Q => 
                           send_ppm1_sig_out_local_count_6_port, QN => n_1007);
   send_ppm1_local_counter1_o_count_reg_7_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N53, C => n129, Q => 
                           send_ppm1_sig_out_local_count_7_port, QN => n_1008);
   send_ppm1_local_counter1_o_count_reg_8_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N54, C => n129, Q => 
                           send_ppm1_sig_out_local_count_8_port, QN => n_1009);
   send_ppm1_local_counter1_o_count_reg_9_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N55, C => n129, Q => 
                           send_ppm1_sig_out_local_count_9_port, QN => n_1010);
   send_ppm1_local_counter1_o_count_reg_10_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N56, C => n129, Q => 
                           send_ppm1_sig_out_local_count_10_port, QN => n_1011)
                           ;
   send_ppm1_local_counter1_o_count_reg_11_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N57, C => n129, Q => 
                           send_ppm1_sig_out_local_count_11_port, QN => n_1012)
                           ;
   send_ppm1_local_counter1_o_count_reg_12_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N58, C => n129, Q => 
                           send_ppm1_sig_out_local_count_12_port, QN => n_1013)
                           ;
   send_ppm1_local_counter1_o_count_reg_13_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N59, C => n129, Q => 
                           send_ppm1_sig_out_local_count_13_port, QN => n_1014)
                           ;
   send_ppm1_local_counter1_o_count_reg_14_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N60, C => n129, Q => 
                           send_ppm1_sig_out_local_count_14_port, QN => n_1015)
                           ;
   send_ppm1_local_counter1_o_count_reg_15_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N61, C => n129, Q => 
                           send_ppm1_sig_out_local_count_15_port, QN => n_1016)
                           ;
   send_ppm1_local_counter1_o_count_reg_16_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N62, C => n129, Q => 
                           send_ppm1_sig_out_local_count_16_port, QN => n_1017)
                           ;
   send_ppm1_local_counter1_o_count_reg_17_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N63, C => n129, Q => 
                           send_ppm1_sig_out_local_count_17_port, QN => n_1018)
                           ;
   send_ppm1_local_counter1_o_count_reg_18_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N64, C => n130, Q => 
                           send_ppm1_sig_out_local_count_18_port, QN => n_1019)
                           ;
   send_ppm1_local_counter1_o_count_reg_19_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N65, C => n129, Q => 
                           send_ppm1_sig_out_local_count_19_port, QN => n_1020)
                           ;
   send_ppm1_local_counter1_v_val_reg_19_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N65, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_19_port, QN => n_1021
                           );
   send_ppm1_local_counter1_v_val_reg_18_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N64, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_18_port, QN => n_1022
                           );
   send_ppm1_local_counter1_v_val_reg_17_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N63, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_17_port, QN => n_1023
                           );
   send_ppm1_local_counter1_v_val_reg_16_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N62, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_16_port, QN => n_1024
                           );
   send_ppm1_local_counter1_v_val_reg_15_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N61, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_15_port, QN => n_1025
                           );
   send_ppm1_local_counter1_v_val_reg_14_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N60, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_14_port, QN => n_1026
                           );
   send_ppm1_local_counter1_v_val_reg_13_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N59, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_13_port, QN => n_1027
                           );
   send_ppm1_local_counter1_v_val_reg_12_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N58, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_12_port, QN => n_1028
                           );
   send_ppm1_local_counter1_v_val_reg_11_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N57, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_11_port, QN => n_1029
                           );
   send_ppm1_local_counter1_v_val_reg_10_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N56, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_10_port, QN => n_1030
                           );
   send_ppm1_local_counter1_v_val_reg_9_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N55, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_9_port, QN => n_1031)
                           ;
   send_ppm1_local_counter1_v_val_reg_8_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N54, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_8_port, QN => n_1032)
                           ;
   send_ppm1_local_counter1_v_val_reg_7_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N53, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_7_port, QN => n_1033)
                           ;
   send_ppm1_local_counter1_v_val_reg_6_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N52, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_6_port, QN => n_1034)
                           ;
   send_ppm1_local_counter1_v_val_reg_5_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N51, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_5_port, QN => n_1035)
                           ;
   send_ppm1_local_counter1_v_val_reg_4_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N50, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_4_port, QN => n_1036)
                           ;
   send_ppm1_local_counter1_v_val_reg_3_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N49, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_3_port, QN => n_1037)
                           ;
   send_ppm1_local_counter1_v_val_reg_2_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N48, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_2_port, QN => n_1038)
                           ;
   send_ppm1_local_counter1_v_val_reg_1_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N47, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_1_port, QN => n_1039)
                           ;
   send_ppm1_local_counter1_v_val_reg_0_inst : DF3 port map( D => 
                           send_ppm1_local_counter1_N46, C => n129, Q => 
                           send_ppm1_local_counter1_v_val_0_port, QN => n_1040)
                           ;
   send_ppm1_sig_reg_storage_reg_13_inst : DFE1 port map( D => sig_reg_14_port,
                           E => n126, C => n130, Q => 
                           send_ppm1_sig_reg_storage_13_port, QN => n_1041);
   send_ppm1_sig_reg_storage_reg_5_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n127, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_5_port, QN => n_1042);
   send_ppm1_sig_reg_storage_reg_6_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n127, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_6_port, QN => n_1043);
   send_ppm1_sig_reg_storage_reg_14_inst : DFE1 port map( D => sig_reg_14_port,
                           E => n126, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_14_port, QN => n_1044);
   send_ppm1_sig_reg_storage_reg_21_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n125, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_21_port, QN => n_1045);
   send_ppm1_sig_reg_storage_reg_22_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n125, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_22_port, QN => n_1046);
   send_ppm1_sig_reg_storage_reg_29_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_29_port, QN => n_1047);
   send_ppm1_sig_reg_storage_reg_30_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_30_port, QN => n_1048);
   send_ppm1_sig_reg_storage_reg_4_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n127, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_4_port, QN => n9);
   send_ppm1_sig_reg_storage_reg_12_inst : DFE1 port map( D => sig_reg_14_port,
                           E => n126, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_12_port, QN => n10);
   send_ppm1_sig_reg_storage_reg_20_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n125, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_20_port, QN => n11);
   send_ppm1_sig_reg_storage_reg_28_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_28_port, QN => n8);
   send_ppm1_sig_reg_storage_reg_2_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n128, C => n130, Q => 
                           send_ppm1_sig_reg_storage_2_port, QN => n_1049);
   send_ppm1_sig_reg_storage_reg_3_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n128, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_3_port, QN => n_1050);
   send_ppm1_sig_reg_storage_reg_10_inst : DFE1 port map( D => sig_reg_14_port,
                           E => n127, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_10_port, QN => n_1051);
   send_ppm1_sig_reg_storage_reg_11_inst : DFE1 port map( D => sig_reg_14_port,
                           E => n126, C => n129, Q => 
                           send_ppm1_sig_reg_storage_11_port, QN => n_1052);
   send_ppm1_sig_reg_storage_reg_18_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n125, C => n129, Q => 
                           send_ppm1_sig_reg_storage_18_port, QN => n_1053);
   send_ppm1_sig_reg_storage_reg_19_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n125, C => n130, Q => 
                           send_ppm1_sig_reg_storage_19_port, QN => n_1054);
   send_ppm1_sig_reg_storage_reg_26_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => n130, Q => 
                           send_ppm1_sig_reg_storage_26_port, QN => n_1055);
   send_ppm1_sig_reg_storage_reg_27_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => n130, Q => 
                           send_ppm1_sig_reg_storage_27_port, QN => n_1056);
   send_ppm1_sig_reg_storage_reg_1_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n128, C => n130, Q => 
                           send_ppm1_sig_reg_storage_1_port, QN => n23);
   send_ppm1_sig_reg_storage_reg_17_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n126, C => n130, Q => 
                           send_ppm1_sig_reg_storage_17_port, QN => n22);
   send_ppm1_sig_reg_storage_reg_9_inst : DFE1 port map( D => sig_reg_14_port, 
                           E => n127, C => n130, Q => 
                           send_ppm1_sig_reg_storage_9_port, QN => n21);
   send_ppm1_sig_reg_storage_reg_25_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n124, C => n130, Q => 
                           send_ppm1_sig_reg_storage_25_port, QN => n20);
   send_ppm1_sig_reg_storage_reg_31_inst : DFE1 port map( D => sig_reg_31_port,
                           E => n124, C => n130, Q => 
                           send_ppm1_sig_reg_storage_31_port, QN => n19);
   send_ppm1_sig_reg_storage_reg_7_inst : DFE1 port map( D => sig_reg_7_port, E
                           => n127, C => n130, Q => 
                           send_ppm1_sig_reg_storage_7_port, QN => n18);
   send_ppm1_sig_reg_storage_reg_23_inst : DFE1 port map( D => i_sel_top(2), E 
                           => n125, C => n130, Q => 
                           send_ppm1_sig_reg_storage_23_port, QN => n17);
   send_ppm1_sig_reg_storage_reg_15_inst : DFE1 port map( D => sig_reg_15_port,
                           E => n126, C => n130, Q => 
                           send_ppm1_sig_reg_storage_15_port, QN => n16);
   send_ppm1_sig_reg_storage_reg_16_inst : DFE1 port map( D => sig_reg_22_port,
                           E => n126, C => n130, Q => 
                           send_ppm1_sig_reg_storage_16_port, QN => n15);
   send_ppm1_sig_reg_storage_reg_8_inst : DFE1 port map( D => sig_reg_14_port, 
                           E => n127, C => n130, Q => 
                           send_ppm1_sig_reg_storage_8_port, QN => n14);
   send_ppm1_sig_reg_storage_reg_24_inst : DFE1 port map( D => sig_reg_30_port,
                           E => n125, C => sig_clk25, Q => 
                           send_ppm1_sig_reg_storage_24_port, QN => n12);
   send_ppm1_sig_reg_storage_reg_0_inst : DFE1 port map( D => sig_reg_6_port, E
                           => n128, C => n130, Q => 
                           send_ppm1_sig_reg_storage_0_port, QN => n13);
   U5 : NOR21 port map( A => n122, B => n25, Q => send_ppm1_local_counter1_N65)
                           ;
   U6 : MUX22 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, B 
                           => n158, S => 
                           send_ppm1_dp_cluster_1_mult_114_A2_8_port, Q => n2);
   U7 : MUX22 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, B 
                           => n178, S => 
                           send_ppm1_dp_cluster_2_mult_117_A2_8_port, Q => n4);
   U8 : MUX22 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, B 
                           => n200, S => 
                           send_ppm1_dp_cluster_4_mult_123_A2_8_port, Q => n5);
   U9 : MUX22 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, B 
                           => n190, S => 
                           send_ppm1_dp_cluster_3_mult_120_A2_8_port, Q => n6);
   U10 : XNR21 port map( A => n151, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, Q 
                           => send_ppm1_dp_cluster_0_N279);
   U11 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, B 
                           => send_ppm1_dp_cluster_0_N279, Q => n56);
   U12 : INV3 port map( A => n54, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port);
   U13 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port, B 
                           => n151, Q => n54);
   U14 : XNR21 port map( A => n151, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, Q 
                           => send_ppm1_dp_cluster_0_N280);
   U15 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, Q 
                           => n151);
   U16 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_12_port, B => n61, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port);
   U17 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, Q 
                           => n61);
   U18 : INV3 port map( A => send_ppm1_dp_cluster_0_N48, Q => n174);
   U19 : INV3 port map( A => n55, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port);
   U20 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, B 
                           => send_ppm1_dp_cluster_0_N280, Q => n55);
   U21 : INV3 port map( A => n53, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_18_port);
   U22 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port, B 
                           => n151, Q => n53);
   U23 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_16_port, Q 
                           => n170);
   U24 : XNR21 port map( A => n151, B => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, Q 
                           => send_ppm1_dp_cluster_0_N281);
   U25 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_15_port, B => n64, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port);
   U26 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, Q 
                           => n64);
   U27 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_13_port, B => n62, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port);
   U28 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, Q 
                           => n62);
   U29 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_14_port, B => n63, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port);
   U30 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, Q 
                           => n63);
   U31 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_11_port, B => n60, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port);
   U32 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, Q 
                           => n60);
   U33 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_12_port, Q => n196);
   U34 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_12_port, B 
                           => n154, Q => send_ppm1_dp_cluster_0_N28);
   U35 : INV3 port map( A => send_ppm1_dp_cluster_0_N45, Q => n180);
   U36 : INV3 port map( A => send_ppm1_dp_cluster_0_N46, Q => n177);
   U37 : INV3 port map( A => send_ppm1_dp_cluster_0_N47, Q => n176);
   U38 : INV3 port map( A => send_ppm1_dp_cluster_0_N49, Q => n173);
   U39 : INV3 port map( A => send_ppm1_dp_cluster_0_N50, Q => n172);
   U40 : INV3 port map( A => send_ppm1_dp_cluster_0_N51, Q => n171);
   U41 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_10_port, B => n28, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port);
   U42 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_12_port, Q => n154);
   U43 : INV3 port map( A => n52, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_17_port);
   U44 : NOR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_16_port, B 
                           => n151, Q => n52);
   U45 : INV3 port map( A => n28, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port);
   U46 : NOR21 port map( A => n160, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, Q 
                           => n28);
   U47 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_2_N250, Q => 
                           send_ppm1_sig_cyclesTrame2_12_port);
   U48 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_3_N235, Q => 
                           send_ppm1_sig_cyclesTrame3_12_port);
   U49 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_1_N265, Q => 
                           send_ppm1_sig_cyclesTrame1_12_port);
   U50 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, 
                           B => send_ppm1_dp_cluster_4_N220, Q => 
                           send_ppm1_sig_cyclesTrame4_12_port);
   U51 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_15_port, B 
                           => n33, Q => send_ppm1_dp_cluster_0_N31);
   U52 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_5_port, B => n59, Q =>
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port);
   U53 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, Q 
                           => n59);
   U54 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_8_port, B => n27, Q =>
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port);
   U55 : NOR21 port map( A => n89, B => n90, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port);
   U56 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port, Q
                           => n89);
   U57 : INV3 port map( A => send_ppm1_dp_cluster_2_N250, Q => n90);
   U58 : NOR21 port map( A => n103, B => n104, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port);
   U59 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port, Q
                           => n103);
   U60 : INV3 port map( A => send_ppm1_dp_cluster_3_N235, Q => n104);
   U61 : NOR21 port map( A => n75, B => n76, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port);
   U62 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port, Q
                           => n75);
   U63 : INV3 port map( A => send_ppm1_dp_cluster_1_N265, Q => n76);
   U64 : NOR21 port map( A => n117, B => n118, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port);
   U65 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port, Q
                           => n117);
   U66 : INV3 port map( A => send_ppm1_dp_cluster_4_N220, Q => n118);
   U67 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_14_port, Q => n194);
   U68 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_14_port, B 
                           => n152, Q => send_ppm1_dp_cluster_0_N30);
   U69 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_10_port, Q => n199);
   U70 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_10_port, B 
                           => n157, Q => send_ppm1_dp_cluster_0_N26);
   U71 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_9_port, Q => n202);
   U72 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_9_port, B 
                           => n160, Q => send_ppm1_dp_cluster_0_N25);
   U73 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_13_port, Q => n195);
   U74 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_13_port, B 
                           => n153, Q => send_ppm1_dp_cluster_0_N29);
   U75 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_11_port, Q => n198);
   U76 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_11_port, B 
                           => n156, Q => send_ppm1_dp_cluster_0_N27);
   U77 : INV3 port map( A => send_ppm1_dp_cluster_0_N41, Q => n184);
   U78 : INV3 port map( A => send_ppm1_dp_cluster_0_N42, Q => n183);
   U79 : INV3 port map( A => send_ppm1_dp_cluster_0_N43, Q => n182);
   U80 : INV3 port map( A => send_ppm1_dp_cluster_0_N44, Q => n181);
   U81 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_9_port, Q => n160);
   U82 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_13_port, Q => n153);
   U83 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_11_port, Q => n156);
   U84 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_14_port, Q => n152);
   U85 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_10_port, Q => n157);
   U86 : INV3 port map( A => n26, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port);
   U87 : NOR21 port map( A => n163, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, Q 
                           => n26);
   U88 : INV3 port map( A => n27, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port);
   U89 : NOR21 port map( A => n162, B => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, Q 
                           => n27);
   U90 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port, 
                           B => send_ppm1_dp_cluster_2_N249, Q => 
                           send_ppm1_sig_cyclesTrame2_13_port);
   U91 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, B
                           => send_ppm1_dp_cluster_2_N253, Q => 
                           send_ppm1_sig_cyclesTrame2_9_port);
   U92 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port, 
                           B => send_ppm1_dp_cluster_2_N251, Q => 
                           send_ppm1_sig_cyclesTrame2_11_port);
   U93 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
                           B => send_ppm1_dp_cluster_3_N234, Q => 
                           send_ppm1_sig_cyclesTrame3_13_port);
   U94 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, B
                           => send_ppm1_dp_cluster_3_N238, Q => 
                           send_ppm1_sig_cyclesTrame3_9_port);
   U95 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port, 
                           B => send_ppm1_dp_cluster_3_N236, Q => 
                           send_ppm1_sig_cyclesTrame3_11_port);
   U96 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port, 
                           B => send_ppm1_dp_cluster_2_N248, Q => 
                           send_ppm1_sig_cyclesTrame2_14_port);
   U97 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port, 
                           B => n4, Q => send_ppm1_sig_cyclesTrame2_10_port);
   U98 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port, 
                           B => send_ppm1_dp_cluster_3_N233, Q => 
                           send_ppm1_sig_cyclesTrame3_14_port);
   U99 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port, 
                           B => n6, Q => send_ppm1_sig_cyclesTrame3_10_port);
   U100 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_1_N268, Q => 
                           send_ppm1_sig_cyclesTrame1_9_port);
   U101 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port,
                           B => send_ppm1_dp_cluster_1_N264, Q => 
                           send_ppm1_sig_cyclesTrame1_13_port);
   U102 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port,
                           B => send_ppm1_dp_cluster_4_N219, Q => 
                           send_ppm1_sig_cyclesTrame4_13_port);
   U103 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, 
                           B => send_ppm1_dp_cluster_4_N223, Q => 
                           send_ppm1_sig_cyclesTrame4_9_port);
   U104 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port,
                           B => send_ppm1_dp_cluster_1_N266, Q => 
                           send_ppm1_sig_cyclesTrame1_11_port);
   U105 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port,
                           B => send_ppm1_dp_cluster_4_N221, Q => 
                           send_ppm1_sig_cyclesTrame4_11_port);
   U106 : XOR21 port map( A => n254, B => n155, Q => 
                           send_ppm1_dp_cluster_1_N265);
   U107 : XOR21 port map( A => n236, B => n197, Q => 
                           send_ppm1_dp_cluster_4_N220);
   U108 : XOR21 port map( A => n248, B => n175, Q => 
                           send_ppm1_dp_cluster_2_N250);
   U109 : XOR21 port map( A => n242, B => n189, Q => 
                           send_ppm1_dp_cluster_3_N235);
   U110 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_1_N263, Q => 
                           send_ppm1_sig_cyclesTrame1_14_port);
   U111 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port,
                           B => send_ppm1_dp_cluster_4_N218, Q => 
                           send_ppm1_sig_cyclesTrame4_14_port);
   U112 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port,
                           B => n2, Q => send_ppm1_sig_cyclesTrame1_10_port);
   U113 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port,
                           B => n5, Q => send_ppm1_sig_cyclesTrame4_10_port);
   U114 : NAND22 port map( A => decoder1_n11, B => n141, Q => sig_reg_14_port);
   U115 : INV3 port map( A => sig_reg_15_port, Q => n141);
   U116 : NOR21 port map( A => n72, B => n73, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port);
   U117 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port, Q
                           => n72);
   U118 : INV3 port map( A => send_ppm1_dp_cluster_1_N268, Q => n73);
   U119 : NOR21 port map( A => n114, B => n115, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port);
   U120 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port, Q
                           => n114);
   U121 : INV3 port map( A => send_ppm1_dp_cluster_4_N223, Q => n115);
   U122 : NOR21 port map( A => n86, B => n87, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port);
   U123 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port, Q
                           => n86);
   U124 : INV3 port map( A => send_ppm1_dp_cluster_2_N253, Q => n87);
   U125 : NOR21 port map( A => n100, B => n101, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port);
   U126 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port, Q
                           => n100);
   U127 : INV3 port map( A => send_ppm1_dp_cluster_3_N238, Q => n101);
   U128 : NOR21 port map( A => n91, B => n92, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port);
   U129 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_13_port, 
                           Q => n91);
   U130 : INV3 port map( A => send_ppm1_dp_cluster_2_N249, Q => n92);
   U131 : NOR21 port map( A => n105, B => n106, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port);
   U132 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_13_port, 
                           Q => n105);
   U133 : INV3 port map( A => send_ppm1_dp_cluster_3_N234, Q => n106);
   U134 : NOR21 port map( A => n77, B => n78, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port);
   U135 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_13_port, 
                           Q => n77);
   U136 : INV3 port map( A => send_ppm1_dp_cluster_1_N264, Q => n78);
   U137 : NOR21 port map( A => n119, B => n120, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port);
   U138 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_13_port, 
                           Q => n119);
   U139 : INV3 port map( A => send_ppm1_dp_cluster_4_N219, Q => n120);
   U140 : NOR21 port map( A => n32, B => n74, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_12_port);
   U141 : INV3 port map( A => send_ppm1_dp_cluster_1_N266, Q => n74);
   U142 : NOR21 port map( A => n47, B => n116, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_12_port);
   U143 : INV3 port map( A => send_ppm1_dp_cluster_4_N221, Q => n116);
   U144 : NOR21 port map( A => n37, B => n88, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_12_port);
   U145 : INV3 port map( A => send_ppm1_dp_cluster_2_N251, Q => n88);
   U146 : NOR21 port map( A => n42, B => n102, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_12_port);
   U147 : INV3 port map( A => send_ppm1_dp_cluster_3_N236, Q => n102);
   U148 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_4_port, B => n58, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port);
   U149 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, Q 
                           => n58);
   U150 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_6_port, Q => n205);
   U151 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_6_port, B 
                           => n163, Q => send_ppm1_dp_cluster_0_N22);
   U152 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_5_port, Q => n206);
   U153 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_5_port, B 
                           => n164, Q => send_ppm1_dp_cluster_0_N21);
   U154 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_7_port, Q => n204);
   U155 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_7_port, B 
                           => n162, Q => send_ppm1_dp_cluster_0_N23);
   U156 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_8_port, Q => n203);
   U157 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_8_port, B 
                           => n161, Q => send_ppm1_dp_cluster_0_N24);
   U158 : INV3 port map( A => send_ppm1_dp_cluster_0_N39, Q => n186);
   U159 : INV3 port map( A => send_ppm1_dp_cluster_0_N40, Q => n185);
   U160 : INV3 port map( A => send_ppm1_N198, Q => n149);
   U161 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_7_port, Q => n162);
   U162 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_8_port, Q => n161);
   U163 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_5_port, Q => n164);
   U164 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_6_port, Q => n163);
   U165 : INV3 port map( A => n38, Q => send_ppm1_sig_cyclesTrame2_15_port);
   U166 : NOR21 port map( A => send_ppm1_dp_cluster_2_N248, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_14_port, Q 
                           => n38);
   U167 : INV3 port map( A => n43, Q => send_ppm1_sig_cyclesTrame3_15_port);
   U168 : NOR21 port map( A => send_ppm1_dp_cluster_3_N233, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_14_port, Q 
                           => n43);
   U169 : INV3 port map( A => n33, Q => send_ppm1_sig_cyclesTrame1_15_port);
   U170 : NOR21 port map( A => send_ppm1_dp_cluster_1_N263, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_14_port, Q 
                           => n33);
   U171 : INV3 port map( A => n48, Q => send_ppm1_sig_cyclesTrame4_15_port);
   U172 : NOR21 port map( A => send_ppm1_dp_cluster_4_N218, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_14_port, Q 
                           => n48);
   U173 : INV3 port map( A => n32, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_11_port);
   U174 : NOR21 port map( A => n2, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_10_port, Q 
                           => n32);
   U175 : INV3 port map( A => n47, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_11_port);
   U176 : NOR21 port map( A => n5, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_10_port, Q 
                           => n47);
   U177 : INV3 port map( A => n37, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_11_port);
   U178 : NOR21 port map( A => n4, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_10_port, Q 
                           => n37);
   U179 : INV3 port map( A => n42, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_11_port);
   U180 : NOR21 port map( A => n6, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_10_port, Q 
                           => n42);
   U181 : BUF2 port map( A => n146, Q => n124);
   U182 : BUF2 port map( A => n146, Q => n125);
   U183 : BUF2 port map( A => n146, Q => n126);
   U184 : BUF2 port map( A => n146, Q => n127);
   U185 : BUF2 port map( A => n146, Q => n128);
   U186 : NOR40 port map( A => n150, B => n283, C => n282, D => n281, Q => 
                           send_ppm1_N198);
   U187 : INV3 port map( A => n269, Q => n150);
   U188 : NAND22 port map( A => n280, B => n279, Q => n281);
   U189 : NAND31 port map( A => n278, B => n277, C => n276, Q => n282);
   U190 : NOR31 port map( A => send_ppm1_n71, B => send_ppm1_n72, C => 
                           send_ppm1_n70, Q => send_ppm1_n69);
   U191 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_8_port);
   U192 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_5_port);
   U193 : XOR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_7_port);
   U194 : NAND31 port map( A => n139, B => n137, C => decoder1_n14, Q => 
                           decoder1_n11);
   U195 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_8_port);
   U196 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_5_port);
   U197 : XOR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_7_port);
   U198 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame2_6_port);
   U199 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame3_6_port);
   U200 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_8_port);
   U201 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_8_port);
   U202 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_5_port);
   U203 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_5_port);
   U204 : XOR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_7_port);
   U205 : XOR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_7_port);
   U206 : NAND41 port map( A => n169, B => n275, C => n274, D => n273, Q => 
                           n283);
   U207 : INV3 port map( A => n270, Q => n169);
   U208 : NOR21 port map( A => n272, B => n271, Q => n273);
   U209 : NAND22 port map( A => n7, B => send_ppm1_N179, Q => n275);
   U210 : XOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_A1_11_port, B =>
                           n247, Q => send_ppm1_dp_cluster_2_N249);
   U211 : NOR21 port map( A => n175, B => n248, Q => n247);
   U212 : XOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_A1_11_port, B =>
                           n241, Q => send_ppm1_dp_cluster_3_N234);
   U213 : NOR21 port map( A => n189, B => n242, Q => n241);
   U214 : XOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_A1_11_port, B =>
                           n253, Q => send_ppm1_dp_cluster_1_N264);
   U215 : NOR21 port map( A => n155, B => n254, Q => n253);
   U216 : XOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_A1_11_port, B =>
                           n235, Q => send_ppm1_dp_cluster_4_N219);
   U217 : NOR21 port map( A => n197, B => n236, Q => n235);
   U218 : XOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_1_N268);
   U219 : XOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_4_N223);
   U220 : XOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_2_N253);
   U221 : XOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, B
                           => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           Q => send_ppm1_dp_cluster_3_N238);
   U222 : XNR21 port map( A => n244, B => 
                           send_ppm1_dp_cluster_2_mult_117_A2_12_port, Q => 
                           send_ppm1_dp_cluster_2_N248);
   U223 : NAND22 port map( A => send_ppm1_dp_cluster_2_mult_117_A1_11_port, B 
                           => n245, Q => n244);
   U224 : NOR21 port map( A => n81, B => n16, Q => 
                           send_ppm1_dp_cluster_2_mult_117_A2_12_port);
   U225 : NOR21 port map( A => n175, B => n246, Q => n245);
   U226 : XNR21 port map( A => n238, B => 
                           send_ppm1_dp_cluster_3_mult_120_A2_12_port, Q => 
                           send_ppm1_dp_cluster_3_N233);
   U227 : NAND22 port map( A => send_ppm1_dp_cluster_3_mult_120_A1_11_port, B 
                           => n239, Q => n238);
   U228 : NOR21 port map( A => n95, B => n17, Q => 
                           send_ppm1_dp_cluster_3_mult_120_A2_12_port);
   U229 : NOR21 port map( A => n189, B => n240, Q => n239);
   U230 : XNR21 port map( A => n250, B => 
                           send_ppm1_dp_cluster_1_mult_114_A2_12_port, Q => 
                           send_ppm1_dp_cluster_1_N263);
   U231 : NAND22 port map( A => send_ppm1_dp_cluster_1_mult_114_A1_11_port, B 
                           => n251, Q => n250);
   U232 : NOR21 port map( A => n67, B => n18, Q => 
                           send_ppm1_dp_cluster_1_mult_114_A2_12_port);
   U233 : NOR21 port map( A => n155, B => n252, Q => n251);
   U234 : XNR21 port map( A => n232, B => 
                           send_ppm1_dp_cluster_4_mult_123_A2_12_port, Q => 
                           send_ppm1_dp_cluster_4_N218);
   U235 : NAND22 port map( A => send_ppm1_dp_cluster_4_mult_123_A1_11_port, B 
                           => n233, Q => n232);
   U236 : NOR21 port map( A => n109, B => n19, Q => 
                           send_ppm1_dp_cluster_4_mult_123_A2_12_port);
   U237 : NOR21 port map( A => n197, B => n234, Q => n233);
   U238 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame1_6_port);
   U239 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, 
                           B => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, 
                           Q => send_ppm1_sig_cyclesTrame4_6_port);
   U240 : XOR21 port map( A => n159, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_1_N266);
   U241 : XOR21 port map( A => n201, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_4_N221);
   U242 : XOR21 port map( A => n179, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_2_N251);
   U243 : XOR21 port map( A => n191, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           send_ppm1_dp_cluster_3_N236);
   U244 : NAND22 port map( A => decoder1_n11, B => n138, Q => sig_reg_6_port);
   U245 : INV3 port map( A => sig_reg_7_port, Q => n138);
   U246 : NAND22 port map( A => decoder1_n11, B => n139, Q => sig_reg_22_port);
   U247 : NAND22 port map( A => decoder1_n11, B => n137, Q => sig_reg_30_port);
   U248 : XNR21 port map( A => send_ppm1_dp_cluster_0_N296, B => n24, Q => 
                           send_ppm1_N179);
   U249 : NOR40 port map( A => n371, B => n370, C => n369, D => n368, Q => 
                           send_ppm1_N148);
   U250 : NAND41 port map( A => n168, B => n355, C => n354, D => n353, Q => 
                           n371);
   U251 : NAND41 port map( A => n359, B => n358, C => n357, D => n356, Q => 
                           n370);
   U252 : NAND41 port map( A => n363, B => n362, C => n361, D => n360, Q => 
                           n369);
   U253 : NOR40 port map( A => n268, B => n267, C => n266, D => n265, Q => n269
                           );
   U254 : NAND22 port map( A => n259, B => n258, Q => n267);
   U255 : NAND22 port map( A => n264, B => n263, Q => n265);
   U256 : NAND31 port map( A => n257, B => n256, C => n255, Q => n268);
   U257 : AOI221 port map( A => n7, B => n3_port, C => n3_port, D => 
                           send_ppm1_N179, Q => n270);
   U258 : NAND22 port map( A => n159, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           n254);
   U259 : NAND22 port map( A => n201, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           n236);
   U260 : NAND22 port map( A => n179, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           n248);
   U261 : NAND22 port map( A => n191, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           n242);
   U262 : INV3 port map( A => send_ppm1_n71, Q => n211);
   U263 : INV3 port map( A => send_ppm1_n60, Q => n146);
   U264 : NOR21 port map( A => n30, B => n68, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port);
   U265 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port, Q 
                           => n68);
   U266 : NOR21 port map( A => n45, B => n110, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port);
   U267 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port, Q 
                           => n110);
   U268 : NOR21 port map( A => n35, B => n82, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port);
   U269 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port, Q 
                           => n82);
   U270 : NOR21 port map( A => n40, B => n96, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port);
   U271 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port, Q 
                           => n96);
   U272 : NOR21 port map( A => n65, B => n66, Q => 
                           send_ppm1_dp_cluster_1_mult_114_A2_8_port);
   U273 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_4_5_port, Q 
                           => n66);
   U274 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_1_port, 
                           Q => n65);
   U275 : NOR21 port map( A => n107, B => n108, Q => 
                           send_ppm1_dp_cluster_4_mult_123_A2_8_port);
   U276 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_4_5_port, Q 
                           => n108);
   U277 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_1_port, 
                           Q => n107);
   U278 : NOR21 port map( A => n79, B => n80, Q => 
                           send_ppm1_dp_cluster_2_mult_117_A2_8_port);
   U279 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_4_5_port, Q 
                           => n80);
   U280 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_1_port, 
                           Q => n79);
   U281 : NOR21 port map( A => n93, B => n94, Q => 
                           send_ppm1_dp_cluster_3_mult_120_A2_8_port);
   U282 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_4_5_port, Q 
                           => n94);
   U283 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_1_port, 
                           Q => n93);
   U284 : NOR21 port map( A => n70, B => n71, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_9_port);
   U285 : INV3 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port, Q
                           => n70);
   U286 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_7_1_port, Q 
                           => n71);
   U287 : NOR21 port map( A => n112, B => n113, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_9_port);
   U288 : INV3 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port, Q
                           => n112);
   U289 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_7_1_port, Q 
                           => n113);
   U290 : NOR21 port map( A => n84, B => n85, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_9_port);
   U291 : INV3 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port, Q
                           => n84);
   U292 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_7_1_port, Q 
                           => n85);
   U293 : NOR21 port map( A => n98, B => n99, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_9_port);
   U294 : INV3 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port, Q
                           => n98);
   U295 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_7_1_port, Q 
                           => n99);
   U296 : NOR21 port map( A => n31, B => n69, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_8_port);
   U297 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_6_1_port, Q 
                           => n69);
   U298 : NOR21 port map( A => n46, B => n111, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_8_port);
   U299 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_6_1_port, Q 
                           => n111);
   U300 : NOR21 port map( A => n36, B => n83, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_8_port);
   U301 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_6_1_port, Q 
                           => n83);
   U302 : NOR21 port map( A => n41, B => n97, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_8_port);
   U303 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_6_1_port, Q 
                           => n97);
   U304 : INV3 port map( A => n50, Q => 
                           send_ppm1_dp_cluster_0_add_3_root_sub_235_cf_carry_2_port);
   U305 : NOR21 port map( A => n15, B => n14, Q => n50);
   U306 : NOR21 port map( A => send_ppm1_sig_cyclesTrame1_3_port, B => n57, Q 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port);
   U307 : INV3 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, Q 
                           => n57);
   U308 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_3_port, Q => n208);
   U309 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port, B 
                           => n166, Q => send_ppm1_dp_cluster_0_N19);
   U310 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_4_port, Q => n207);
   U311 : XOR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_4_port, B 
                           => n165, Q => send_ppm1_dp_cluster_0_N20);
   U312 : INV3 port map( A => n51, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_2_port);
   U313 : INV3 port map( A => send_ppm1_dp_cluster_0_N38, Q => n187);
   U314 : NOR21 port map( A => n24, B => send_ppm1_dp_cluster_0_N296, Q => n51)
                           ;
   U315 : NAND22 port map( A => n179, B => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_6_5_port, Q => 
                           n246);
   U316 : NAND22 port map( A => n191, B => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_6_5_port, Q => 
                           n240);
   U317 : NAND22 port map( A => n159, B => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_6_5_port, Q => 
                           n252);
   U318 : NAND22 port map( A => n201, B => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_6_5_port, Q => 
                           n234);
   U319 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_7_5_port, Q 
                           => n175);
   U320 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_7_5_port, Q 
                           => n189);
   U321 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_7_5_port, Q 
                           => n155);
   U322 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_7_5_port, Q 
                           => n197);
   U323 : NOR21 port map( A => n7, B => n15, Q => n306);
   U324 : NOR21 port map( A => n7, B => n14, Q => n328);
   U325 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n122);
   U326 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n121);
   U327 : NAND22 port map( A => decoder1_n8, B => decoder1_n12, Q => 
                           sig_reg_15_port);
   U328 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_2_port, Q => n167);
   U329 : NOR21 port map( A => n7, B => n12, Q => n284);
   U330 : INV3 port map( A => send_ppm1_n72, Q => n145);
   U331 : INV3 port map( A => send_ppm1_n76, Q => n148);
   U332 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_3_port, Q => n166);
   U333 : INV3 port map( A => send_ppm1_sig_cyclesTrame1_4_port, Q => n165);
   U334 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, Q 
                           => n158);
   U335 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, Q 
                           => n200);
   U336 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, Q 
                           => n178);
   U337 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, Q 
                           => n190);
   U338 : INV3 port map( A => n249, Q => n159);
   U339 : NAND22 port map( A => send_ppm1_dp_cluster_1_mult_114_A2_8_port, B =>
                           send_ppm1_dp_cluster_1_mult_114_SUMB_5_5_port, Q => 
                           n249);
   U340 : INV3 port map( A => n231, Q => n201);
   U341 : NAND22 port map( A => send_ppm1_dp_cluster_4_mult_123_A2_8_port, B =>
                           send_ppm1_dp_cluster_4_mult_123_SUMB_5_5_port, Q => 
                           n231);
   U342 : INV3 port map( A => n243, Q => n179);
   U343 : NAND22 port map( A => send_ppm1_dp_cluster_2_mult_117_A2_8_port, B =>
                           send_ppm1_dp_cluster_2_mult_117_SUMB_5_5_port, Q => 
                           n243);
   U344 : INV3 port map( A => n237, Q => n191);
   U345 : NAND22 port map( A => send_ppm1_dp_cluster_3_mult_120_A2_8_port, B =>
                           send_ppm1_dp_cluster_3_mult_120_SUMB_5_5_port, Q => 
                           n237);
   U346 : BUF2 port map( A => send_ppm1_local_counter1_n22, Q => n123);
   U347 : XOR21 port map( A => n14, B => n15, Q => n24);
   U348 : INV3 port map( A => n31, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_7_port);
   U349 : NOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_1_sub_114_cf_carry_6_port, Q
                           => n31);
   U350 : INV3 port map( A => n46, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_7_port);
   U351 : NOR21 port map( A => send_ppm1_dp_cluster_4_mult_123_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_4_sub_123_cf_carry_6_port, Q
                           => n46);
   U352 : INV3 port map( A => n36, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_7_port);
   U353 : NOR21 port map( A => send_ppm1_dp_cluster_2_mult_117_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_2_sub_117_cf_carry_6_port, Q
                           => n36);
   U354 : INV3 port map( A => n41, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_7_port);
   U355 : NOR21 port map( A => send_ppm1_dp_cluster_3_mult_120_SUMB_5_1_port, B
                           => send_ppm1_dp_cluster_3_sub_120_cf_carry_6_port, Q
                           => n41);
   U356 : INV3 port map( A => send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, 
                           Q => n81);
   U357 : INV3 port map( A => send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, 
                           Q => n95);
   U358 : INV3 port map( A => send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, 
                           Q => n67);
   U359 : INV3 port map( A => send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, 
                           Q => n109);
   U360 : NOR21 port map( A => n122, B => n214, Q => 
                           send_ppm1_local_counter1_N63);
   U361 : INV3 port map( A => send_ppm1_local_counter1_N23, Q => n214);
   U362 : NOR21 port map( A => n122, B => n216, Q => 
                           send_ppm1_local_counter1_N61);
   U363 : INV3 port map( A => send_ppm1_local_counter1_N21, Q => n216);
   U364 : NOR21 port map( A => n122, B => n218, Q => 
                           send_ppm1_local_counter1_N59);
   U365 : INV3 port map( A => send_ppm1_local_counter1_N19, Q => n218);
   U366 : NOR21 port map( A => n122, B => n220, Q => 
                           send_ppm1_local_counter1_N57);
   U367 : INV3 port map( A => send_ppm1_local_counter1_N17, Q => n220);
   U368 : NOR21 port map( A => n122, B => n222, Q => 
                           send_ppm1_local_counter1_N55);
   U369 : INV3 port map( A => send_ppm1_local_counter1_N15, Q => n222);
   U370 : NOR21 port map( A => n122, B => n224, Q => 
                           send_ppm1_local_counter1_N53);
   U371 : INV3 port map( A => send_ppm1_local_counter1_N13, Q => n224);
   U372 : NOR21 port map( A => n121, B => n225, Q => 
                           send_ppm1_local_counter1_N52);
   U373 : INV3 port map( A => send_ppm1_local_counter1_N12, Q => n225);
   U374 : NOR21 port map( A => n121, B => n226, Q => 
                           send_ppm1_local_counter1_N51);
   U375 : INV3 port map( A => send_ppm1_local_counter1_N11, Q => n226);
   U376 : NOR21 port map( A => n121, B => n227, Q => 
                           send_ppm1_local_counter1_N50);
   U377 : INV3 port map( A => send_ppm1_local_counter1_N10, Q => n227);
   U378 : NOR21 port map( A => n121, B => n228, Q => 
                           send_ppm1_local_counter1_N49);
   U379 : INV3 port map( A => send_ppm1_local_counter1_N9, Q => n228);
   U380 : NOR21 port map( A => n121, B => n229, Q => 
                           send_ppm1_local_counter1_N48);
   U381 : INV3 port map( A => send_ppm1_local_counter1_N8, Q => n229);
   U382 : NOR21 port map( A => n121, B => n230, Q => 
                           send_ppm1_local_counter1_N47);
   U383 : INV3 port map( A => send_ppm1_local_counter1_N7, Q => n230);
   U384 : NOR21 port map( A => n123, B => n213, Q => 
                           send_ppm1_local_counter1_N64);
   U385 : INV3 port map( A => send_ppm1_local_counter1_N24, Q => n213);
   U386 : NOR21 port map( A => n123, B => n215, Q => 
                           send_ppm1_local_counter1_N62);
   U387 : INV3 port map( A => send_ppm1_local_counter1_N22_port, Q => n215);
   U388 : NOR21 port map( A => n123, B => n217, Q => 
                           send_ppm1_local_counter1_N60);
   U389 : INV3 port map( A => send_ppm1_local_counter1_N20, Q => n217);
   U390 : NOR21 port map( A => n123, B => n219, Q => 
                           send_ppm1_local_counter1_N58);
   U391 : INV3 port map( A => send_ppm1_local_counter1_N18, Q => n219);
   U392 : NOR21 port map( A => n123, B => n221, Q => 
                           send_ppm1_local_counter1_N56);
   U393 : INV3 port map( A => send_ppm1_local_counter1_N16, Q => n221);
   U394 : NOR21 port map( A => n123, B => n223, Q => 
                           send_ppm1_local_counter1_N54);
   U395 : INV3 port map( A => send_ppm1_local_counter1_N14, Q => n223);
   U396 : INV3 port map( A => send_ppm1_n70, Q => n135);
   U397 : INV3 port map( A => n350, Q => n168);
   U398 : NOR21 port map( A => n7, B => n13, Q => n350);
   U399 : BUF6 port map( A => sig_clk25, Q => n129);
   U400 : NOR21 port map( A => n129, B => n131, Q => N3);
   U401 : INV3 port map( A => i_reset_n_top, Q => n131);
   U402 : NAND41 port map( A => send_ppm1_n82, B => send_ppm1_n83, C => 
                           send_ppm1_n84, D => send_ppm1_n85, Q => 
                           send_ppm1_n71);
   U403 : NOR21 port map( A => send_ppm1_sig_out_local_count_16_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => 
                           send_ppm1_n82);
   U404 : NOR31 port map( A => send_ppm1_n86, B => send_ppm1_n87, C => 
                           send_ppm1_n88, Q => send_ppm1_n85);
   U405 : NOR31 port map( A => send_ppm1_sig_out_local_count_17_port, B => 
                           send_ppm1_sig_out_local_count_19_port, C => 
                           send_ppm1_sig_out_local_count_18_port, Q => 
                           send_ppm1_n83);
   U406 : XOR21 port map( A => send_ppm1_sig_reg_storage_8_port, B => 
                           send_ppm1_sig_reg_storage_9_port, Q => 
                           send_ppm1_sig_cyclesTrame2_2_port);
   U407 : NOR31 port map( A => send_ppm1_sig_state_0_port, B => 
                           send_ppm1_sig_state_1_port, C => send_ppm1_n57, Q =>
                           send_ppm1_n72);
   U408 : XOR21 port map( A => send_ppm1_sig_reg_storage_16_port, B => 
                           send_ppm1_sig_reg_storage_17_port, Q => 
                           send_ppm1_sig_cyclesTrame3_2_port);
   U409 : NOR31 port map( A => send_ppm1_current_state_0_port, B => 
                           send_ppm1_current_state_2_port, C => send_ppm1_n53, 
                           Q => send_ppm1_n76);
   U410 : OAI2111 port map( A => n142, B => decoder1_n10, C => decoder1_n13, D 
                           => decoder1_n12, Q => sig_reg_7_port);
   U411 : INV3 port map( A => decoder1_n14, Q => n142);
   U412 : NAND22 port map( A => i_sel_top(2), B => decoder1_n14, Q => 
                           decoder1_n13);
   U413 : NAND41 port map( A => n342, B => n345, C => n344, D => n343, Q => 
                           n346);
   U414 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n343);
   U415 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n345);
   U416 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n344);
   U417 : NAND41 port map( A => n320, B => n323, C => n322, D => n321, Q => 
                           n324);
   U418 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n321);
   U419 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n323);
   U420 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n322);
   U421 : NAND41 port map( A => n364, B => n367, C => n366, D => n365, Q => 
                           n368);
   U422 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n365);
   U423 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n367);
   U424 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n366);
   U425 : NAND41 port map( A => n298, B => n301, C => n300, D => n299, Q => 
                           n302);
   U426 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_13_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n299);
   U427 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_15_port, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n301);
   U428 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_14_port, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n300);
   U429 : NOR40 port map( A => send_ppm1_sig_out_local_count_5_port, B => n212,
                           C => send_ppm1_sig_out_local_count_4_port, D => 
                           send_ppm1_sig_out_local_count_2_port, Q => 
                           send_ppm1_n84);
   U430 : INV3 port map( A => send_ppm1_n90, Q => n212);
   U431 : NOR21 port map( A => send_ppm1_sig_out_local_count_9_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => 
                           send_ppm1_n90);
   U432 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_10_port, Q => 
                           send_ppm1_sig_cyclesTrame2_3_port);
   U433 : XNR21 port map( A => send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_11_port, Q => 
                           send_ppm1_sig_cyclesTrame2_4_port);
   U434 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n342);
   U435 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n320);
   U436 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n364);
   U437 : NOR40 port map( A => send_ppm1_sig_out_local_count_19_port, B => 
                           send_ppm1_sig_out_local_count_18_port, C => 
                           send_ppm1_sig_out_local_count_17_port, D => 
                           send_ppm1_sig_out_local_count_16_port, Q => n298);
   U438 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_18_port, Q => 
                           send_ppm1_sig_cyclesTrame3_3_port);
   U439 : XNR21 port map( A => send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_19_port, Q => 
                           send_ppm1_sig_cyclesTrame3_4_port);
   U440 : INV3 port map( A => send_ppm1_N169, Q => n193);
   U441 : AOI311 port map( A => send_ppm1_N148, B => send_ppm1_n58, C => 
                           send_ppm1_sig_state_0_port, D => send_ppm1_n92, Q =>
                           send_ppm1_n91);
   U442 : NOR40 port map( A => n305, B => n304, C => n303, D => n302, Q => 
                           send_ppm1_N169);
   U443 : NAND41 port map( A => n341, B => n340, C => n339, D => n338, Q => 
                           n347);
   U444 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n338);
   U445 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n339);
   U446 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n340);
   U447 : NAND41 port map( A => n319, B => n318, C => n317, D => n316, Q => 
                           n325);
   U448 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n316);
   U449 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n317);
   U450 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n318);
   U451 : NAND41 port map( A => n297, B => n296, C => n295, D => n294, Q => 
                           n303);
   U452 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n294);
   U453 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n295);
   U454 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n296);
   U455 : NAND41 port map( A => send_ppm1_sig_out_local_count_11_port, B => 
                           send_ppm1_sig_out_local_count_10_port, C => 
                           send_ppm1_n89, D => 
                           send_ppm1_sig_out_local_count_0_port, Q => 
                           send_ppm1_n86);
   U456 : NOR21 port map( A => send_ppm1_sig_out_local_count_14_port, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => 
                           send_ppm1_n89);
   U457 : XOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => 
                           send_ppm1_sig_reg_storage_25_port, Q => 
                           send_ppm1_sig_cyclesTrame4_2_port);
   U458 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => 
                           send_ppm1_sig_reg_storage_1_port, Q => 
                           send_ppm1_sig_cyclesTrame1_2_port);
   U459 : NAND41 port map( A => n337, B => n336, C => n335, D => n334, Q => 
                           n348);
   U460 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n334);
   U461 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n336);
   U462 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n335);
   U463 : NAND41 port map( A => n315, B => n314, C => n313, D => n312, Q => 
                           n326);
   U464 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n312);
   U465 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n314);
   U466 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n313);
   U467 : NAND41 port map( A => n293, B => n292, C => n291, D => n290, Q => 
                           n304);
   U468 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n290);
   U469 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n292);
   U470 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n291);
   U471 : XOR21 port map( A => send_ppm1_sig_reg_storage_4_port, B => 
                           send_ppm1_sig_reg_storage_0_port, Q => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_4_1_port);
   U472 : XOR21 port map( A => send_ppm1_sig_reg_storage_28_port, B => 
                           send_ppm1_sig_reg_storage_24_port, Q => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_4_1_port);
   U473 : XOR21 port map( A => send_ppm1_sig_reg_storage_12_port, B => 
                           send_ppm1_sig_reg_storage_8_port, Q => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_4_1_port);
   U474 : XOR21 port map( A => send_ppm1_sig_reg_storage_20_port, B => 
                           send_ppm1_sig_reg_storage_16_port, Q => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_4_1_port);
   U475 : XNR21 port map( A => n13, B => send_ppm1_sig_reg_storage_24_port, Q 
                           => send_ppm1_dp_cluster_0_N296);
   U476 : NAND41 port map( A => n188, B => n333, C => n332, D => n331, Q => 
                           n349);
   U477 : INV3 port map( A => n328, Q => n188);
   U478 : NOR21 port map( A => n330, B => n329, Q => n331);
   U479 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n332);
   U480 : NAND41 port map( A => n192, B => n311, C => n310, D => n309, Q => 
                           n327);
   U481 : INV3 port map( A => n306, Q => n192);
   U482 : NOR21 port map( A => n308, B => n307, Q => n309);
   U483 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n310);
   U484 : NAND41 port map( A => n210, B => n289, C => n288, D => n287, Q => 
                           n305);
   U485 : INV3 port map( A => n284, Q => n210);
   U486 : NOR21 port map( A => n286, B => n285, Q => n287);
   U487 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n288);
   U488 : XOR21 port map( A => send_ppm1_sig_reg_storage_15_port, B => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_2_mult_117_A1_11_port);
   U489 : XOR21 port map( A => send_ppm1_sig_reg_storage_23_port, B => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_3_mult_120_A1_11_port);
   U490 : XOR21 port map( A => send_ppm1_sig_reg_storage_7_port, B => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_1_mult_114_A1_11_port);
   U491 : XOR21 port map( A => send_ppm1_sig_reg_storage_31_port, B => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_7_5_port, Q 
                           => send_ppm1_dp_cluster_4_mult_123_A1_11_port);
   U492 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_2_port, Q => 
                           send_ppm1_sig_cyclesTrame1_3_port);
   U493 : XNR21 port map( A => send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_3_port, Q => 
                           send_ppm1_sig_cyclesTrame1_4_port);
   U494 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, 
                           B => send_ppm1_sig_reg_storage_26_port, Q => 
                           send_ppm1_sig_cyclesTrame4_3_port);
   U495 : XNR21 port map( A => send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, 
                           B => send_ppm1_sig_reg_storage_27_port, Q => 
                           send_ppm1_sig_cyclesTrame4_4_port);
   U496 : AOI221 port map( A => send_ppm1_n63, B => 
                           send_ppm1_current_state_1_port, C => send_ppm1_n62, 
                           D => send_ppm1_current_state_2_port, Q => 
                           send_ppm1_n60);
   U497 : NOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => n13, Q 
                           => n49);
   U498 : NAND22 port map( A => i_reset_n_top, B => send_ppm1_n79, Q => 
                           send_ppm1_n70);
   U499 : NOR21 port map( A => n147, B => send_ppm1_current_state_2_port, Q => 
                           send_ppm1_n79);
   U500 : INV3 port map( A => send_ppm1_n62, Q => n147);
   U501 : OAI2111 port map( A => n137, B => decoder1_n8, C => decoder1_n9, D =>
                           decoder1_n10, Q => sig_reg_31_port);
   U502 : NAND22 port map( A => i_sel_top(3), B => n140, Q => decoder1_n9);
   U503 : INV3 port map( A => i_sel_top(1), Q => n140);
   U504 : OAI2111 port map( A => send_ppm1_N198, B => n148, C => send_ppm1_n78,
                           D => i_reset_n_top, Q => send_ppm1_N82_port);
   U505 : NAND31 port map( A => send_ppm1_n72, B => n211, C => send_ppm1_n79, Q
                           => send_ppm1_n78);
   U506 : OAI2111 port map( A => send_ppm1_n64, B => send_ppm1_n80, C => 
                           send_ppm1_n81, D => i_reset_n_top, Q => 
                           send_ppm1_N81_port);
   U507 : NAND22 port map( A => send_ppm1_n63, B => send_ppm1_n53, Q => 
                           send_ppm1_n80);
   U508 : NAND31 port map( A => n211, B => n145, C => send_ppm1_n79, Q => 
                           send_ppm1_n81);
   U509 : NOR21 port map( A => send_ppm1_n55, B => 
                           send_ppm1_current_state_2_port, Q => send_ppm1_n63);
   U510 : NOR21 port map( A => n143, B => i_sel_top(1), Q => decoder1_n14);
   U511 : NAND31 port map( A => n262, B => n261, C => n260, Q => n266);
   U512 : XNR21 port map( A => send_ppm1_N193, B => 
                           send_ppm1_sig_out_local_count_15_port, Q => n262);
   U513 : XNR21 port map( A => send_ppm1_N192, B => 
                           send_ppm1_sig_out_local_count_14_port, Q => n261);
   U514 : XNR21 port map( A => send_ppm1_N194, B => 
                           send_ppm1_sig_out_local_count_16_port, Q => n260);
   U515 : XOR21 port map( A => send_ppm1_sig_cyclesTrame2_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n330);
   U516 : NAND31 port map( A => send_ppm1_sig_out_local_count_1_port, B => 
                           send_ppm1_sig_out_local_count_12_port, C => 
                           send_ppm1_sig_out_local_count_3_port, Q => 
                           send_ppm1_n87);
   U517 : XOR21 port map( A => send_ppm1_sig_cyclesTrame3_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n308);
   U518 : XOR21 port map( A => send_ppm1_sig_cyclesTrame4_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n286);
   U519 : XOR21 port map( A => send_ppm1_N180, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n272);
   U520 : XOR21 port map( A => send_ppm1_sig_cyclesTrame2_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n329);
   U521 : XOR21 port map( A => send_ppm1_sig_cyclesTrame3_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n307);
   U522 : XOR21 port map( A => send_ppm1_sig_cyclesTrame4_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n285);
   U523 : XOR21 port map( A => send_ppm1_N181, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n271);
   U524 : INV3 port map( A => send_ppm1_n66, Q => n132);
   U525 : INV3 port map( A => send_ppm1_n69, Q => n136);
   U526 : NAND22 port map( A => send_ppm1_sig_state_0_port, B => send_ppm1_n58,
                           Q => send_ppm1_n65);
   U527 : NOR21 port map( A => n12, B => n20, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port);
   U528 : NOR21 port map( A => n13, B => n23, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port);
   U529 : NOR21 port map( A => n12, B => n20, Q => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_1_5_port);
   U530 : NOR21 port map( A => n13, B => n23, Q => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_1_5_port);
   U531 : NOR21 port map( A => n8, B => n12, Q => 
                           send_ppm1_dp_cluster_4_mult_123_CARRYB_4_1_port);
   U532 : XOR21 port map( A => send_ppm1_sig_reg_storage_24_port, B => 
                           send_ppm1_sig_reg_storage_25_port, Q => 
                           send_ppm1_dp_cluster_4_mult_123_SUMB_1_5_port);
   U533 : NOR21 port map( A => n9, B => n13, Q => 
                           send_ppm1_dp_cluster_1_mult_114_CARRYB_4_1_port);
   U534 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => 
                           send_ppm1_sig_reg_storage_1_port, Q => 
                           send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port);
   U535 : NOR21 port map( A => n14, B => n21, Q => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_1_5_port);
   U536 : NOR21 port map( A => n15, B => n22, Q => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_1_5_port);
   U537 : NOR21 port map( A => n10, B => n14, Q => 
                           send_ppm1_dp_cluster_2_mult_117_CARRYB_4_1_port);
   U538 : XOR21 port map( A => send_ppm1_sig_reg_storage_8_port, B => 
                           send_ppm1_sig_reg_storage_9_port, Q => 
                           send_ppm1_dp_cluster_2_mult_117_SUMB_1_5_port);
   U539 : NOR21 port map( A => n11, B => n15, Q => 
                           send_ppm1_dp_cluster_3_mult_120_CARRYB_4_1_port);
   U540 : XOR21 port map( A => send_ppm1_sig_reg_storage_16_port, B => 
                           send_ppm1_sig_reg_storage_17_port, Q => 
                           send_ppm1_dp_cluster_3_mult_120_SUMB_1_5_port);
   U541 : NOR21 port map( A => send_ppm1_current_state_0_port, B => 
                           send_ppm1_current_state_1_port, Q => send_ppm1_n62);
   U542 : NOR21 port map( A => n14, B => n21, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port);
   U543 : NOR21 port map( A => n15, B => n22, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port);
   U544 : NOR21 port map( A => send_ppm1_dp_cluster_1_mult_114_SUMB_1_5_port, B
                           => n13, Q => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_3_port);
   U545 : XNR21 port map( A => send_ppm1_N185, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n279);
   U546 : XNR21 port map( A => send_ppm1_N195, B => 
                           send_ppm1_sig_out_local_count_17_port, Q => n263);
   U547 : XNR21 port map( A => send_ppm1_dp_cluster_0_N280, B => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_17_port, Q 
                           => send_ppm1_N195);
   U548 : XNR21 port map( A => send_ppm1_N190, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n258);
   U549 : XNR21 port map( A => send_ppm1_N184, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n276);
   U550 : XNR21 port map( A => send_ppm1_N189, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n255);
   U551 : NAND22 port map( A => send_ppm1_sig_out_local_count_8_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => 
                           send_ppm1_n88);
   U552 : AOI211 port map( A => n135, B => send_ppm1_n58, C => send_ppm1_n66, Q
                           => send_ppm1_n67);
   U553 : NAND41 port map( A => send_ppm1_n69, B => send_ppm1_sig_state_1_port,
                           C => send_ppm1_sig_state_0_port, D => send_ppm1_n57,
                           Q => send_ppm1_n68);
   U554 : INV3 port map( A => n49, Q => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_2_port);
   U555 : INV3 port map( A => send_ppm1_sig_cyclesTrame4_2_port, Q => n209);
   U556 : XOR21 port map( A => send_ppm1_sig_reg_storage_0_port, B => n167, Q 
                           => send_ppm1_dp_cluster_0_N18);
   U557 : NAND22 port map( A => i_sel_top(1), B => i_sel_top(0), Q => 
                           decoder1_n12);
   U558 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n337);
   U559 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n315);
   U560 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n359);
   U561 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_8_port, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n293);
   U562 : XNR21 port map( A => send_ppm1_sig_cyclesTrame2_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n341);
   U563 : XNR21 port map( A => send_ppm1_sig_cyclesTrame3_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n319);
   U564 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n363);
   U565 : XNR21 port map( A => send_ppm1_sig_cyclesTrame4_12_port, B => 
                           send_ppm1_sig_out_local_count_12_port, Q => n297);
   U566 : XNR21 port map( A => send_ppm1_N191, B => 
                           send_ppm1_sig_out_local_count_13_port, Q => n259);
   U567 : XNR21 port map( A => send_ppm1_N186, B => 
                           send_ppm1_sig_out_local_count_8_port, Q => n280);
   U568 : XNR21 port map( A => send_ppm1_N196, B => 
                           send_ppm1_sig_out_local_count_18_port, Q => n264);
   U569 : XNR21 port map( A => send_ppm1_dp_cluster_0_N279, B => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_18_port, Q 
                           => send_ppm1_N196);
   U570 : NAND22 port map( A => i_sel_top(3), B => n139, Q => decoder1_n10);
   U571 : XNR21 port map( A => send_ppm1_N187, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n256);
   U572 : XNR21 port map( A => send_ppm1_N182, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n277);
   U573 : NAND22 port map( A => i_sel_top(1), B => n143, Q => decoder1_n8);
   U574 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_6_port, B => 
                           send_ppm1_sig_out_local_count_6_port, Q => n357);
   U575 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_7_port, B => 
                           send_ppm1_sig_out_local_count_7_port, Q => n358);
   U576 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_2_port, B => 
                           send_ppm1_sig_out_local_count_2_port, Q => n354);
   U577 : XNR21 port map( A => send_ppm1_N183, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n278);
   U578 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_11_port, B => 
                           send_ppm1_sig_out_local_count_11_port, Q => n362);
   U579 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_10_port, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n361);
   U580 : XNR21 port map( A => send_ppm1_N188, B => 
                           send_ppm1_sig_out_local_count_10_port, Q => n257);
   U581 : XNR21 port map( A => send_ppm1_N197, B => 
                           send_ppm1_sig_out_local_count_19_port, Q => n274);
   U582 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port, B 
                           => send_ppm1_dp_cluster_0_N278, Q => send_ppm1_N197)
                           ;
   U583 : INV3 port map( A => n56, Q => 
                           send_ppm1_dp_cluster_0_sub_0_root_sub_235_cf_carry_19_port);
   U584 : XNR21 port map( A => 
                           send_ppm1_dp_cluster_0_add_1_root_sub_235_cf_carry_19_port, B 
                           => 
                           send_ppm1_dp_cluster_0_sub_4_root_sub_235_cf_carry_16_port, Q 
                           => send_ppm1_dp_cluster_0_N278);
   U585 : NAND22 port map( A => i_reset_n_top, B => n144, Q => 
                           send_ppm1_local_counter1_n22);
   U586 : INV3 port map( A => send_ppm1_sig_in_init, Q => n144);
   U587 : OAI2111 port map( A => n148, B => n149, C => send_ppm1_n60, D => 
                           send_ppm1_n61, Q => send_ppm1_sig_in_init);
   U588 : AOI221 port map( A => n211, B => send_ppm1_n62, C => send_ppm1_n63, D
                           => send_ppm1_n64, Q => send_ppm1_n61);
   U589 : INV3 port map( A => n44, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port);
   U590 : NOR21 port map( A => send_ppm1_sig_reg_storage_26_port, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_3_port, Q =>
                           n44);
   U591 : INV3 port map( A => n34, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port);
   U592 : NOR21 port map( A => send_ppm1_sig_reg_storage_10_port, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_3_port, Q =>
                           n34);
   U593 : INV3 port map( A => n39, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port);
   U594 : NOR21 port map( A => send_ppm1_sig_reg_storage_18_port, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_3_port, Q =>
                           n39);
   U595 : INV3 port map( A => n29, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port);
   U596 : NOR21 port map( A => send_ppm1_sig_reg_storage_2_port, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_3_port, Q =>
                           n29);
   U597 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_9_port, B => 
                           send_ppm1_sig_out_local_count_9_port, Q => n360);
   U598 : XNR21 port map( A => send_ppm1_sig_cyclesTrame1_5_port, B => 
                           send_ppm1_sig_out_local_count_5_port, Q => n356);
   U599 : INV3 port map( A => n30, Q => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_5_port);
   U600 : NOR21 port map( A => send_ppm1_sig_reg_storage_3_port, B => 
                           send_ppm1_dp_cluster_1_sub_114_cf_carry_4_port, Q =>
                           n30);
   U601 : INV3 port map( A => n45, Q => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_5_port);
   U602 : NOR21 port map( A => send_ppm1_sig_reg_storage_27_port, B => 
                           send_ppm1_dp_cluster_4_sub_123_cf_carry_4_port, Q =>
                           n45);
   U603 : INV3 port map( A => n35, Q => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_5_port);
   U604 : NOR21 port map( A => send_ppm1_sig_reg_storage_11_port, B => 
                           send_ppm1_dp_cluster_2_sub_117_cf_carry_4_port, Q =>
                           n35);
   U605 : INV3 port map( A => n40, Q => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_5_port);
   U606 : NOR21 port map( A => send_ppm1_sig_reg_storage_19_port, B => 
                           send_ppm1_dp_cluster_3_sub_120_cf_carry_4_port, Q =>
                           n40);
   U607 : INV3 port map( A => i_sel_top(2), Q => n139);
   U608 : NOR21 port map( A => send_ppm1_n93, B => send_ppm1_n58, Q => 
                           send_ppm1_n92);
   U609 : AOI221 port map( A => send_ppm1_N156, B => send_ppm1_n59, C => 
                           send_ppm1_N163, D => send_ppm1_sig_state_0_port, Q 
                           => send_ppm1_n93);
   U610 : NOR40 port map( A => n327, B => n326, C => n325, D => n324, Q => 
                           send_ppm1_N163);
   U611 : NOR40 port map( A => n349, B => n348, C => n347, D => n346, Q => 
                           send_ppm1_N156);
   U612 : INV3 port map( A => i_sel_top(3), Q => n137);
   U613 : NOR21 port map( A => n121, B => send_ppm1_local_counter1_v_val_0_port
                           , Q => send_ppm1_local_counter1_N46);
   U614 : NOR21 port map( A => n352, B => n351, Q => n353);
   U615 : XOR21 port map( A => send_ppm1_sig_cyclesTrame1_4_port, B => 
                           send_ppm1_sig_out_local_count_4_port, Q => n351);
   U616 : XOR21 port map( A => send_ppm1_sig_cyclesTrame1_3_port, B => 
                           send_ppm1_sig_out_local_count_3_port, Q => n352);
   U617 : INV3 port map( A => send_ppm1_n73, Q => n133);
   U618 : OAI2111 port map( A => n211, B => send_ppm1_n70, C => send_ppm1_n74, 
                           D => send_ppm1_n75, Q => send_ppm1_n73);
   U619 : NAND31 port map( A => send_ppm1_n76, B => n149, C => i_reset_n_top, Q
                           => send_ppm1_n74);
   U620 : NAND31 port map( A => send_ppm1_n63, B => send_ppm1_n53, C => 
                           i_reset_n_top, Q => send_ppm1_n75);
   U621 : XNR21 port map( A => send_ppm1_local_counter1_add_34_carry_19_port, B
                           => send_ppm1_local_counter1_v_val_19_port, Q => n25)
                           ;
   U622 : INV3 port map( A => i_sel_top(0), Q => n143);
   U623 : INV3 port map( A => send_ppm1_n77, Q => n134);
   U624 : NAND31 port map( A => i_reset_n_top, B => send_ppm1_n76, C => 
                           send_ppm1_N198, Q => send_ppm1_n77);
   U625 : BUF2 port map( A => sig_clk25, Q => n130);
   U626 : OAI222 port map( A => n3_port, B => n7, C => n12, D => n3_port, Q => 
                           n289);
   U627 : OAI222 port map( A => n3_port, B => n7, C => n15, D => n3_port, Q => 
                           n311);
   U628 : OAI222 port map( A => n3_port, B => n7, C => n14, D => n3_port, Q => 
                           n333);
   U629 : OAI222 port map( A => n3_port, B => n7, C => n13, D => n3_port, Q => 
                           n355);

end SYN_rtl;
